// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.8.0.115.3
// Netlist written on Thu Apr 06 15:21:53 2017
//
// Verilog Description of module SPI_loopback_Top
//

module SPI_loopback_Top (CS, SCK, MOSI, MISO, HALL_A_OUT, HALL_B_OUT, 
            HALL_C_OUT, LED1, LED2, LED3, LED4, clkout, H_A_m1, 
            H_B_m1, H_C_m1, MA_m1, MB_m1, MC_m1, H_A_m2, H_B_m2, 
            H_C_m2, MA_m2, MB_m2, MC_m2, H_A_m3, H_B_m3, H_C_m3, 
            MA_m3, MB_m3, MC_m3, H_A_m4, H_B_m4, H_C_m4, MA_m4, 
            MB_m4, MC_m4);   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(24[8:24])
    input CS;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(27[2:4])
    input SCK;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(28[2:5])
    input MOSI;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(29[2:6])
    output MISO;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(30[2:6])
    output HALL_A_OUT;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(33[2:12])
    output HALL_B_OUT;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(34[2:12])
    output HALL_C_OUT;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(35[2:12])
    output LED1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(38[2:6])
    output LED2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(39[2:6])
    output LED3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(40[2:6])
    output LED4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(41[2:6])
    output clkout;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    input H_A_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(47[2:8])
    input H_B_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(48[2:8])
    input H_C_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(49[2:8])
    output [1:0]MA_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(50[2:7])
    output [1:0]MB_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(51[2:7])
    output [1:0]MC_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(52[2:7])
    input H_A_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(55[2:8])
    input H_B_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(56[2:8])
    input H_C_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(57[2:8])
    output [1:0]MA_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(58[2:7])
    output [1:0]MB_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(59[2:7])
    output [1:0]MC_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(60[2:7])
    input H_A_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(63[2:8])
    input H_B_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(64[2:8])
    input H_C_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(65[2:8])
    output [1:0]MA_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(66[2:7])
    output [1:0]MB_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(67[2:7])
    output [1:0]MC_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(68[2:7])
    input H_A_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(71[2:8])
    input H_B_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(72[2:8])
    input H_C_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(73[2:8])
    output [1:0]MA_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(74[2:7])
    output [1:0]MB_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(75[2:7])
    output [1:0]MC_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(76[2:7])
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(88[9:16])
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(30[4:14])
    
    wire GND_net, VCC_net, HALL_A_OUT_c_c, HALL_B_OUT_c_c, HALL_C_OUT_c_c, 
        LED1_c, LED2_c, LED3_c, LED4_c, H_A_m1_c, H_B_m1_c, H_C_m1_c, 
        MA_m1_c_1, MA_m1_c_0, MB_m1_c_1, MB_m1_c_0, MC_m1_c_1, MC_m1_c_0, 
        H_A_m2_c, H_B_m2_c, H_C_m2_c, MA_m2_c_1, MA_m2_c_0, MB_m2_c_1, 
        MB_m2_c_0, MC_m2_c_1, MC_m2_c_0, H_A_m3_c, H_B_m3_c, H_C_m3_c, 
        MA_m3_c_1, MA_m3_c_0, MB_m3_c_1, MB_m3_c_0, MC_m3_c_1, MC_m3_c_0, 
        H_A_m4_c, H_B_m4_c, H_C_m4_c, MA_m4_c_1, MA_m4_c_0, MB_m4_c_1, 
        MB_m4_c_0, MC_m4_c_1, MC_m4_c_0, rst, enable_m1, enable_m2, 
        enable_m3, enable_m4;
    wire [20:0]speed_set_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(99[9:21])
    wire [20:0]speed_set_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(100[9:21])
    wire [20:0]speed_set_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(101[9:21])
    wire [20:0]speed_set_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(102[9:21])
    wire [20:0]speed_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(104[9:17])
    wire [20:0]speed_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(105[9:17])
    wire [20:0]speed_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(106[9:17])
    wire [20:0]speed_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(107[9:17])
    wire [2:0]hallsense_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(110[9:21])
    wire [2:0]hallsense_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(111[9:21])
    wire [2:0]hallsense_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(112[9:21])
    wire [2:0]hallsense_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(113[9:21])
    
    wire PWM_m1, PWM_m2, PWM_m3, PWM_m4;
    wire [9:0]PWMdut_m1;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(120[9:18])
    wire [9:0]PWMdut_m2;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(121[9:18])
    wire [9:0]PWMdut_m3;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(122[9:18])
    wire [9:0]PWMdut_m4;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(123[9:18])
    
    wire dir_m1, dir_m2, dir_m3, dir_m4;
    wire [13:0]start_cnt;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(135[9:18])
    
    wire free_m1, free_m2, free_m3, free_m4;
    wire [95:0]send_buffer;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(67[10:21])
    
    wire n3082, n3140, n3058, n3046, n9, n3010, n2952, n20053, 
        n2928, n2916, n2964, n4216, n2880, n2822, n4215, n2798, 
        n2786, n20586, n20051;
    wire [95:0]send_buffer_95__N_346;
    
    wire MISO_N_624, n4213, n4209, n4193, n4182, n3176;
    wire [28:0]intgOut3;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(70[9:17])
    wire [28:0]backOut2;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(79[9:17])
    wire [28:0]backOut3;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(80[9:17])
    
    wire n4184, n4185, n4186, n4187, n4189, n4190, n4191, n4192, 
        n4219, n4220;
    wire [25:0]subOut_24__N_1135;
    
    wire n4201, n4218, n4183, n4188, n4214, n20537, n21, n19, 
        n13, n19704, n13_adj_1939, n13_adj_1940, n18847, n20525, 
        n18846, n18845, n18844, n18843, n18842, n18841, n20041, 
        n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4202, 
        n4203, n4204, n4208, n4210, n4211, n4212, n4227, n19062, 
        n4226, n4225, n18995, n4224, n4223, n4133, n19061, n2834, 
        n22, n4222, n4229, n3094, n4228, n3188, n3212, n3270, 
        n3224, n19454, n4217, n4221, n4884, n6, n20030, n62, 
        n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
        n73, n74, n75, n10082, clkout_c_enable_219, n19700, n21_adj_1941, 
        n19_adj_1942, clkout_c_enable_257, n3, n13_adj_1943, n19702, 
        n21_adj_1944, n19_adj_1945, n34, n30, n32, n5, n31, n7, 
        n14, n13_adj_1946, n10, n13_adj_1947, n10_adj_1948, n13_adj_1949, 
        n10_adj_1950, n19_adj_1951, n13_adj_1952, n10_adj_1953, n13_adj_1954, 
        n10_adj_1955, n19698, n13_adj_1956, n21920, n21918, n21917, 
        n21_adj_1957, n21913, n19_adj_1958, n21911, clkout_c_enable_244, 
        n21910, n19706, n21908, n21907, n21906, n21_adj_1959, n21905, 
        n21902, n21900, n21899, n22378, n22383, n21865, n21864, 
        n21857, n21851, n21837, n21835;
    
    VHI i2 (.Z(VCC_net));
    OSCH OSCInst0 (.STDBY(GND_net), .OSC(clkout_c)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCInst0.NOM_FREQ = "38.00";
    OB MA_m2_pad_0 (.I(MA_m2_c_0), .O(MA_m2[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(58[2:7])
    LUT4 mux_2095_i2_3_lut (.A(n4203), .B(n4228), .C(n19454), .Z(subOut_24__N_1135[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i2_3_lut.init = 16'hacac;
    LUT4 mux_2095_i3_3_lut (.A(n4202), .B(n4227), .C(n19454), .Z(subOut_24__N_1135[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i3_3_lut.init = 16'hacac;
    LUT4 mux_2095_i4_3_lut (.A(n4201), .B(n4226), .C(n19454), .Z(subOut_24__N_1135[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i4_3_lut.init = 16'hacac;
    LUT4 mux_2095_i5_3_lut (.A(n4200), .B(n4225), .C(n19454), .Z(subOut_24__N_1135[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i5_3_lut.init = 16'hacac;
    LUT4 mux_2095_i6_3_lut (.A(n4199), .B(n4224), .C(n19454), .Z(subOut_24__N_1135[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i6_3_lut.init = 16'hacac;
    LUT4 mux_2095_i7_3_lut (.A(n4198), .B(n4223), .C(n19454), .Z(subOut_24__N_1135[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i7_3_lut.init = 16'hacac;
    LUT4 mux_2095_i8_3_lut (.A(n4197), .B(n4222), .C(n19454), .Z(subOut_24__N_1135[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i8_3_lut.init = 16'hacac;
    LUT4 i2269_4_lut_rep_417 (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18995), .Z(n21837)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2269_4_lut_rep_417.init = 16'hccc8;
    LUT4 mux_2095_i9_3_lut (.A(n4196), .B(n4221), .C(n19454), .Z(subOut_24__N_1135[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i9_3_lut.init = 16'hacac;
    LUT4 i8961_1_lut_4_lut (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18995), .Z(clkout_c_enable_257)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i8961_1_lut_4_lut.init = 16'h3337;
    LUT4 mux_2095_i10_3_lut (.A(n4195), .B(n4220), .C(n19454), .Z(subOut_24__N_1135[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i10_3_lut.init = 16'hacac;
    LUT4 mux_2095_i11_3_lut (.A(n4194), .B(n4219), .C(n19454), .Z(subOut_24__N_1135[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i11_3_lut.init = 16'hacac;
    LUT4 mux_2095_i12_3_lut (.A(n4193), .B(n4218), .C(n19454), .Z(subOut_24__N_1135[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i12_3_lut.init = 16'hacac;
    LUT4 mux_2095_i13_3_lut (.A(n4192), .B(n4217), .C(n19454), .Z(subOut_24__N_1135[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i13_3_lut.init = 16'hacac;
    LUT4 mux_2095_i14_3_lut (.A(n4191), .B(n4216), .C(n19454), .Z(subOut_24__N_1135[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i14_3_lut.init = 16'hacac;
    LUT4 mux_2095_i15_3_lut (.A(n4190), .B(n4215), .C(n19454), .Z(subOut_24__N_1135[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i15_3_lut.init = 16'hacac;
    LUT4 mux_2095_i16_3_lut (.A(n4189), .B(n4214), .C(n19454), .Z(subOut_24__N_1135[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i16_3_lut.init = 16'hacac;
    LUT4 mux_2095_i17_3_lut (.A(n4188), .B(n4213), .C(n19454), .Z(subOut_24__N_1135[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i17_3_lut.init = 16'hacac;
    LUT4 mux_2095_i18_3_lut (.A(n4187), .B(n4212), .C(n19454), .Z(subOut_24__N_1135[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i18_3_lut.init = 16'hacac;
    LUT4 mux_2095_i19_3_lut (.A(n4186), .B(n4211), .C(n19454), .Z(subOut_24__N_1135[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i19_3_lut.init = 16'hacac;
    LUT4 mux_2095_i20_3_lut (.A(n4185), .B(n4210), .C(n19454), .Z(subOut_24__N_1135[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i20_3_lut.init = 16'hacac;
    OB HALL_B_OUT_pad (.I(HALL_B_OUT_c_c), .O(HALL_B_OUT));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(34[2:12])
    OB HALL_A_OUT_pad (.I(HALL_A_OUT_c_c), .O(HALL_A_OUT));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(33[2:12])
    OB MA_m2_pad_1 (.I(MA_m2_c_1), .O(MA_m2[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(58[2:7])
    IB H_B_m1_pad (.I(H_B_m1), .O(H_B_m1_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(48[2:8])
    LUT4 mux_2095_i21_3_lut (.A(n4184), .B(n4209), .C(n19454), .Z(subOut_24__N_1135[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i21_3_lut.init = 16'hacac;
    OBZ n4883_pad (.I(MISO_N_624), .T(n4884), .O(MISO));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(64[1] 216[13])
    IB H_A_m1_pad (.I(H_A_m1), .O(H_A_m1_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(47[2:8])
    IB HALL_C_OUT_c_pad (.I(MOSI), .O(HALL_C_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(29[2:6])
    IB HALL_B_OUT_c_pad (.I(SCK), .O(HALL_B_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(28[2:5])
    IB HALL_A_OUT_c_pad (.I(CS), .O(HALL_A_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(27[2:4])
    OB MC_m4_pad_0 (.I(MC_m4_c_0), .O(MC_m4[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(76[2:7])
    LUT4 mux_2095_i22_3_lut (.A(n4183), .B(n4208), .C(n19454), .Z(subOut_24__N_1135[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i22_3_lut.init = 16'hacac;
    OB MC_m4_pad_1 (.I(MC_m4_c_1), .O(MC_m4[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(76[2:7])
    OB MB_m4_pad_0 (.I(MB_m4_c_0), .O(MB_m4[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(75[2:7])
    LUT4 mux_2095_i25_3_lut (.A(n4182), .B(n4208), .C(n19454), .Z(subOut_24__N_1135[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i25_3_lut.init = 16'hacac;
    OB MB_m4_pad_1 (.I(MB_m4_c_1), .O(MB_m4[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(75[2:7])
    OB MC_m1_pad_0 (.I(MC_m1_c_0), .O(MC_m1[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(52[2:7])
    OB MC_m1_pad_1 (.I(MC_m1_c_1), .O(MC_m1[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(52[2:7])
    OB MA_m4_pad_0 (.I(MA_m4_c_0), .O(MA_m4[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_0 (.I(MB_m1_c_0), .O(MB_m1[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(51[2:7])
    OB MA_m4_pad_1 (.I(MA_m4_c_1), .O(MA_m4[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_1 (.I(MB_m1_c_1), .O(MB_m1[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(51[2:7])
    OB MC_m3_pad_0 (.I(MC_m3_c_0), .O(MC_m3[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(68[2:7])
    IB H_C_m4_pad (.I(H_C_m4), .O(H_C_m4_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(73[2:8])
    OB MA_m1_pad_0 (.I(MA_m1_c_0), .O(MA_m1[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(50[2:7])
    OB MC_m3_pad_1 (.I(MC_m3_c_1), .O(MC_m3[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(68[2:7])
    IB H_B_m4_pad (.I(H_B_m4), .O(H_B_m4_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(72[2:8])
    OB MA_m1_pad_1 (.I(MA_m1_c_1), .O(MA_m1[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(50[2:7])
    OB MB_m3_pad_0 (.I(MB_m3_c_0), .O(MB_m3[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(67[2:7])
    IB H_A_m4_pad (.I(H_A_m4), .O(H_A_m4_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(71[2:8])
    OB clkout_pad (.I(clkout_c), .O(clkout));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    OB MB_m3_pad_1 (.I(MB_m3_c_1), .O(MB_m3[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(67[2:7])
    IB H_C_m3_pad (.I(H_C_m3), .O(H_C_m3_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(65[2:8])
    OB LED4_pad (.I(LED4_c), .O(LED4));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(41[2:6])
    OB MA_m3_pad_0 (.I(MA_m3_c_0), .O(MA_m3[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(66[2:7])
    IB H_B_m3_pad (.I(H_B_m3), .O(H_B_m3_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(64[2:8])
    OB LED3_pad (.I(LED3_c), .O(LED3));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(40[2:6])
    OB MA_m3_pad_1 (.I(MA_m3_c_1), .O(MA_m3[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(66[2:7])
    IB H_A_m3_pad (.I(H_A_m3), .O(H_A_m3_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(63[2:8])
    OB LED2_pad (.I(LED2_c), .O(LED2));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(39[2:6])
    OB MC_m2_pad_0 (.I(MC_m2_c_0), .O(MC_m2[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(60[2:7])
    IB H_C_m2_pad (.I(H_C_m2), .O(H_C_m2_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(57[2:8])
    OB LED1_pad (.I(LED1_c), .O(LED1));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(38[2:6])
    OB MC_m2_pad_1 (.I(MC_m2_c_1), .O(MC_m2[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(60[2:7])
    IB H_B_m2_pad (.I(H_B_m2), .O(H_B_m2_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(56[2:8])
    OB HALL_C_OUT_pad (.I(HALL_C_OUT_c_c), .O(HALL_C_OUT));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(35[2:12])
    OB MB_m2_pad_0 (.I(MB_m2_c_0), .O(MB_m2[0]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(59[2:7])
    IB H_A_m2_pad (.I(H_A_m2), .O(H_A_m2_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(55[2:8])
    OB MB_m2_pad_1 (.I(MB_m2_c_1), .O(MB_m2[1]));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(59[2:7])
    IB H_C_m1_pad (.I(H_C_m1), .O(H_C_m1_c));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(49[2:8])
    FD1P3AX start_cnt_2059__i0 (.D(n75), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i0.GSR = "DISABLED";
    LUT4 m1_lut (.Z(n22378)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    CLKDIV CLKDIV_I (.clkout_c(clkout_c), .clk_1mhz(clk_1mhz), .pwm_clk(pwm_clk), 
           .GND_net(GND_net), .clk_N_683(clk_N_683));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(288[14:20])
    LUT4 i1_2_lut_4_lut (.A(send_buffer[94]), .B(speed_m1[19]), .C(n21864), 
         .D(n21865), .Z(send_buffer_95__N_346[94])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(73[10:15])
    defparam i1_2_lut_4_lut.init = 16'h00ca;
    FD1S3AX rst_13_rep_513 (.D(n21837), .CK(clkout_c), .Q(clkout_c_enable_244));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_13_rep_513.GSR = "DISABLED";
    LUT4 i13178_4_lut (.A(n4133), .B(speed_m3[19]), .C(n21857), .D(speed_m4[19]), 
         .Z(n3)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i13178_4_lut.init = 16'hcac0;
    COMMUTATION_U8 COM_I_M1 (.MB_m1_c_0(MB_m1_c_0), .clkout_c(clkout_c), 
            .MC_m1_c_0(MC_m1_c_0), .MA_m1_c_0(MA_m1_c_0), .LED1_c(LED1_c), 
            .MA_m1_c_1(MA_m1_c_1), .n20053(n20053), .n2880(n2880), .MC_m1_c_1(MC_m1_c_1), 
            .n2834(n2834), .n2822(n2822), .MB_m1_c_1(MB_m1_c_1), .n2798(n2798), 
            .n2786(n2786), .enable_m1(enable_m1), .n21920(n21920), .PWM_m1(PWM_m1), 
            .n21918(n21918), .n21917(n21917), .free_m1(free_m1));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(305[13:24])
    LUT4 i40_4_lut (.A(backOut2[0]), .B(n9), .C(n21851), .D(backOut3[0]), 
         .Z(n22)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i40_4_lut.init = 16'h3a0a;
    LUT4 i28_4_lut (.A(backOut2[5]), .B(n9), .C(n21851), .D(backOut3[5]), 
         .Z(n13_adj_1946)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i28_4_lut.init = 16'h3a0a;
    LUT4 i28_4_lut_adj_201 (.A(backOut2[4]), .B(n9), .C(n21851), .D(backOut3[4]), 
         .Z(n13_adj_1947)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i28_4_lut_adj_201.init = 16'h3a0a;
    LUT4 i28_4_lut_adj_202 (.A(backOut2[3]), .B(n9), .C(n21851), .D(backOut3[3]), 
         .Z(n13_adj_1949)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i28_4_lut_adj_202.init = 16'h3a0a;
    LUT4 i28_4_lut_adj_203 (.A(backOut2[2]), .B(n9), .C(n21851), .D(backOut3[2]), 
         .Z(n13_adj_1952)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i28_4_lut_adj_203.init = 16'h3a0a;
    LUT4 i28_4_lut_adj_204 (.A(backOut2[1]), .B(n9), .C(n21851), .D(backOut3[1]), 
         .Z(n13_adj_1954)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i28_4_lut_adj_204.init = 16'h3a0a;
    FD1S3AX rst_13_rep_512 (.D(n21837), .CK(clkout_c), .Q(clkout_c_enable_219));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_13_rep_512.GSR = "DISABLED";
    COMMUTATION_U7 COM_I_M2 (.MB_m2_c_0(MB_m2_c_0), .clkout_c(clkout_c), 
            .MC_m2_c_0(MC_m2_c_0), .MA_m2_c_0(MA_m2_c_0), .LED2_c(LED2_c), 
            .MA_m2_c_1(MA_m2_c_1), .n20041(n20041), .n3010(n3010), .MC_m2_c_1(MC_m2_c_1), 
            .n2964(n2964), .n2952(n2952), .MB_m2_c_1(MB_m2_c_1), .n2928(n2928), 
            .n2916(n2916), .enable_m2(enable_m2), .n21913(n21913), .PWM_m2(PWM_m2), 
            .n21911(n21911), .n21910(n21910), .free_m2(free_m2));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(315[13:24])
    COMMUTATION_U6 COM_I_M3 (.MB_m3_c_0(MB_m3_c_0), .clkout_c(clkout_c), 
            .MC_m3_c_0(MC_m3_c_0), .MA_m3_c_0(MA_m3_c_0), .LED3_c(LED3_c), 
            .MA_m3_c_1(MA_m3_c_1), .n20051(n20051), .n3140(n3140), .MC_m3_c_1(MC_m3_c_1), 
            .n3094(n3094), .n3082(n3082), .MB_m3_c_1(MB_m3_c_1), .n3058(n3058), 
            .n3046(n3046), .enable_m3(enable_m3), .n21908(n21908), .PWM_m3(PWM_m3), 
            .n21906(n21906), .n21905(n21905), .free_m3(free_m3));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(325[13:24])
    FD1S3AX rst_13_rep_511 (.D(n21837), .CK(clkout_c), .Q(n22383));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_13_rep_511.GSR = "DISABLED";
    FD1S3AX rst_13 (.D(n21837), .CK(clkout_c), .Q(rst));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_13.GSR = "DISABLED";
    GSR GSR_INST (.GSR(n22383));
    LUT4 mux_2095_i1_3_lut (.A(n4204), .B(n4229), .C(n19454), .Z(subOut_24__N_1135[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam mux_2095_i1_3_lut.init = 16'hacac;
    LUT4 i3_4_lut (.A(n19062), .B(start_cnt[10]), .C(start_cnt[9]), .D(start_cnt[8]), 
         .Z(n18995)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_205 (.A(n19061), .B(n6), .C(start_cnt[6]), .D(start_cnt[4]), 
         .Z(n19062)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_205.init = 16'hfefc;
    L6MUX21 i18 (.D0(n34), .D1(n31), .SD(n20537), .Z(n14));
    L6MUX21 i17 (.D0(n19706), .D1(n19), .SD(n20537), .Z(n13));
    LUT4 i3_4_lut_adj_206 (.A(start_cnt[0]), .B(start_cnt[3]), .C(start_cnt[2]), 
         .D(start_cnt[1]), .Z(n19061)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_206.init = 16'hfffe;
    L6MUX21 i17_adj_207 (.D0(n19704), .D1(n19_adj_1958), .SD(n20537), 
            .Z(n13_adj_1940));
    LUT4 i2_2_lut (.A(start_cnt[7]), .B(start_cnt[5]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    L6MUX21 i17_adj_208 (.D0(n19702), .D1(n19_adj_1951), .SD(n20537), 
            .Z(n13_adj_1956));
    L6MUX21 i17_adj_209 (.D0(n19700), .D1(n19_adj_1945), .SD(n20537), 
            .Z(n13_adj_1943));
    L6MUX21 i17_adj_210 (.D0(n19698), .D1(n19_adj_1942), .SD(n20537), 
            .Z(n13_adj_1939));
    PFUMX i13182 (.BLUT(n3), .ALUT(n5), .C0(n20586), .Z(n7));
    CCU2D start_cnt_2059_add_4_15 (.A0(start_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18847), .S0(n62));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_15.INIT0 = 16'hfaaa;
    defparam start_cnt_2059_add_4_15.INIT1 = 16'h0000;
    defparam start_cnt_2059_add_4_15.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_15.INJECT1_1 = "NO";
    CCU2D start_cnt_2059_add_4_13 (.A0(start_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18846), .COUT(n18847), .S0(n64), .S1(n63));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_13.INIT0 = 16'hfaaa;
    defparam start_cnt_2059_add_4_13.INIT1 = 16'hfaaa;
    defparam start_cnt_2059_add_4_13.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_13.INJECT1_1 = "NO";
    CCU2D start_cnt_2059_add_4_11 (.A0(start_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18845), .COUT(n18846), .S0(n66), .S1(n65));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_11.INIT0 = 16'hfaaa;
    defparam start_cnt_2059_add_4_11.INIT1 = 16'hfaaa;
    defparam start_cnt_2059_add_4_11.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_11.INJECT1_1 = "NO";
    CCU2D start_cnt_2059_add_4_9 (.A0(start_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18844), .COUT(n18845), .S0(n68), .S1(n67));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_9.INIT0 = 16'hfaaa;
    defparam start_cnt_2059_add_4_9.INIT1 = 16'hfaaa;
    defparam start_cnt_2059_add_4_9.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_9.INJECT1_1 = "NO";
    CCU2D start_cnt_2059_add_4_7 (.A0(start_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18843), .COUT(n18844), .S0(n70), .S1(n69));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_7.INIT0 = 16'hfaaa;
    defparam start_cnt_2059_add_4_7.INIT1 = 16'hfaaa;
    defparam start_cnt_2059_add_4_7.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_7.INJECT1_1 = "NO";
    CCU2D start_cnt_2059_add_4_5 (.A0(start_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18842), .COUT(n18843), .S0(n72), .S1(n71));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_5.INIT0 = 16'hfaaa;
    defparam start_cnt_2059_add_4_5.INIT1 = 16'hfaaa;
    defparam start_cnt_2059_add_4_5.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_5.INJECT1_1 = "NO";
    PFUMX i49 (.BLUT(n22), .ALUT(n30), .C0(n20525), .Z(n31));
    PFUMX i37 (.BLUT(n13_adj_1946), .ALUT(n21), .C0(n20525), .Z(n19));
    PFUMX i37_adj_211 (.BLUT(n13_adj_1947), .ALUT(n21_adj_1957), .C0(n20525), 
          .Z(n19_adj_1958));
    PFUMX i37_adj_212 (.BLUT(n13_adj_1949), .ALUT(n21_adj_1959), .C0(n20525), 
          .Z(n19_adj_1951));
    CCU2D start_cnt_2059_add_4_3 (.A0(start_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18841), .COUT(n18842), .S0(n74), .S1(n73));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_3.INIT0 = 16'hfaaa;
    defparam start_cnt_2059_add_4_3.INIT1 = 16'hfaaa;
    defparam start_cnt_2059_add_4_3.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_3.INJECT1_1 = "NO";
    PFUMX i37_adj_213 (.BLUT(n13_adj_1952), .ALUT(n21_adj_1944), .C0(n20525), 
          .Z(n19_adj_1945));
    PFUMX i37_adj_214 (.BLUT(n13_adj_1954), .ALUT(n21_adj_1941), .C0(n20525), 
          .Z(n19_adj_1942));
    LUT4 i1746_3_lut_rep_479 (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .Z(n21899)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(128[9:15])
    defparam i1746_3_lut_rep_479.init = 16'h4242;
    LUT4 i18393_2_lut_4_lut (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .D(free_m4), .Z(n3270)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(128[9:15])
    defparam i18393_2_lut_4_lut.init = 16'hffbd;
    CCU2D start_cnt_2059_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18841), .S1(n75));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059_add_4_1.INIT0 = 16'hF000;
    defparam start_cnt_2059_add_4_1.INIT1 = 16'h0555;
    defparam start_cnt_2059_add_4_1.INJECT1_0 = "NO";
    defparam start_cnt_2059_add_4_1.INJECT1_1 = "NO";
    COMMUTATION COM_I_M4 (.MB_m4_c_0(MB_m4_c_0), .clkout_c(clkout_c), .MC_m4_c_0(MC_m4_c_0), 
            .MA_m4_c_0(MA_m4_c_0), .LED4_c(LED4_c), .MA_m4_c_1(MA_m4_c_1), 
            .n20030(n20030), .n3270(n3270), .MC_m4_c_1(MC_m4_c_1), .n3224(n3224), 
            .n3212(n3212), .MB_m4_c_1(MB_m4_c_1), .n3188(n3188), .n3176(n3176), 
            .enable_m4(enable_m4), .n21902(n21902), .PWM_m4(PWM_m4), .n21900(n21900), 
            .n21899(n21899), .free_m4(free_m4));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(335[13:24])
    LUT4 i1654_3_lut_rep_485 (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .Z(n21905)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(127[9:15])
    defparam i1654_3_lut_rep_485.init = 16'h4242;
    LUT4 i18376_2_lut_4_lut (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .D(free_m3), .Z(n3140)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(127[9:15])
    defparam i18376_2_lut_4_lut.init = 16'hffbd;
    LUT4 i1562_3_lut_rep_490 (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .Z(n21910)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(126[9:15])
    defparam i1562_3_lut_rep_490.init = 16'h4242;
    LUT4 i18395_2_lut_4_lut (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .D(free_m2), .Z(n3010)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(126[9:15])
    defparam i18395_2_lut_4_lut.init = 16'hffbd;
    LUT4 i7784_2_lut (.A(n21837), .B(n62), .Z(n10082)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam i7784_2_lut.init = 16'heeee;
    PFUMX i52 (.BLUT(n32), .ALUT(intgOut3[0]), .C0(n21835), .Z(n34));
    PFUMX i27 (.BLUT(n10_adj_1955), .ALUT(intgOut3[1]), .C0(n21835), .Z(n19698));
    PFUMX i27_adj_215 (.BLUT(n10_adj_1953), .ALUT(intgOut3[2]), .C0(n21835), 
          .Z(n19700));
    PFUMX i27_adj_216 (.BLUT(n10_adj_1950), .ALUT(intgOut3[3]), .C0(n21835), 
          .Z(n19702));
    PFUMX i27_adj_217 (.BLUT(n10_adj_1948), .ALUT(intgOut3[4]), .C0(n21835), 
          .Z(n19704));
    PFUMX i27_adj_218 (.BLUT(n10), .ALUT(intgOut3[5]), .C0(n21835), .Z(n19706));
    HALL_U3 HALL_I_M3 (.clk_1mhz(clk_1mhz), .\speed_m3[0] (speed_m3[0]), 
            .hallsense_m3({hallsense_m3}), .clkout_c_enable_244(clkout_c_enable_244), 
            .H_A_m3_c(H_A_m3_c), .H_B_m3_c(H_B_m3_c), .H_C_m3_c(H_C_m3_c), 
            .clkout_c_enable_219(clkout_c_enable_219), .\speed_m3[1] (speed_m3[1]), 
            .\speed_m3[2] (speed_m3[2]), .\speed_m3[3] (speed_m3[3]), .\speed_m3[4] (speed_m3[4]), 
            .\speed_m3[5] (speed_m3[5]), .\speed_m3[6] (speed_m3[6]), .\speed_m3[7] (speed_m3[7]), 
            .\speed_m3[8] (speed_m3[8]), .\speed_m3[9] (speed_m3[9]), .\speed_m3[10] (speed_m3[10]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_m3[12] (speed_m3[12]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_m3[14] (speed_m3[14]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_m3[16] (speed_m3[16]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_m3[18] (speed_m3[18]), 
            .\speed_m3[19] (speed_m3[19]), .n22378(n22378), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(322[14:18])
    LUT4 i1470_3_lut_rep_497 (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .Z(n21917)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(125[9:15])
    defparam i1470_3_lut_rep_497.init = 16'h4242;
    LUT4 i18397_2_lut_4_lut (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .D(free_m1), .Z(n2880)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(125[9:15])
    defparam i18397_2_lut_4_lut.init = 16'hffbd;
    PWMGENERATOR PWM_I_M4 (.PWM_m4(PWM_m4), .pwm_clk(pwm_clk), .free_m4(free_m4), 
            .clkout_c_enable_244(clkout_c_enable_244), .PWMdut_m4({PWMdut_m4}), 
            .GND_net(GND_net), .hallsense_m4({hallsense_m4}), .n21900(n21900), 
            .enable_m4(enable_m4), .n3224(n3224), .n21902(n21902), .n3188(n3188));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(338[13:25])
    PWMGENERATOR_U0 PWM_I_M3 (.PWM_m3(PWM_m3), .pwm_clk(pwm_clk), .free_m3(free_m3), 
            .clkout_c_enable_219(clkout_c_enable_219), .PWMdut_m3({PWMdut_m3}), 
            .GND_net(GND_net), .hallsense_m3({hallsense_m3}), .n21906(n21906), 
            .enable_m3(enable_m3), .n3094(n3094), .n21907(n21907), .n20051(n20051), 
            .n21908(n21908), .n3058(n3058));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(328[13:25])
    HALL_U5 HALL_I_M1 (.clk_1mhz(clk_1mhz), .\speed_m1[0] (speed_m1[0]), 
            .hallsense_m1({hallsense_m1}), .clkout_c_enable_219(clkout_c_enable_219), 
            .clkout_c_enable_244(clkout_c_enable_244), .H_A_m1_c(H_A_m1_c), 
            .H_B_m1_c(H_B_m1_c), .H_C_m1_c(H_C_m1_c), .\speed_m1[1] (speed_m1[1]), 
            .\speed_m1[2] (speed_m1[2]), .\speed_m1[3] (speed_m1[3]), .\speed_m1[4] (speed_m1[4]), 
            .\speed_m1[5] (speed_m1[5]), .\speed_m1[6] (speed_m1[6]), .\speed_m1[7] (speed_m1[7]), 
            .\speed_m1[8] (speed_m1[8]), .\speed_m1[9] (speed_m1[9]), .\speed_m1[10] (speed_m1[10]), 
            .\speed_m1[11] (speed_m1[11]), .\speed_m1[12] (speed_m1[12]), 
            .\speed_m1[13] (speed_m1[13]), .\speed_m1[14] (speed_m1[14]), 
            .\speed_m1[15] (speed_m1[15]), .\speed_m1[16] (speed_m1[16]), 
            .\speed_m1[17] (speed_m1[17]), .\speed_m1[18] (speed_m1[18]), 
            .\speed_m1[19] (speed_m1[19]), .n22378(n22378), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(302[14:18])
    PWMGENERATOR_U1 PWM_I_M2 (.GND_net(GND_net), .PWM_m2(PWM_m2), .pwm_clk(pwm_clk), 
            .free_m2(free_m2), .clkout_c_enable_219(clkout_c_enable_219), 
            .PWMdut_m2({PWMdut_m2}), .hallsense_m2({hallsense_m2}), .n21911(n21911), 
            .enable_m2(enable_m2), .n2964(n2964), .n21913(n21913), .n2928(n2928));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(318[13:25])
    PWMGENERATOR_U2 PWM_I_M1 (.GND_net(GND_net), .PWM_m1(PWM_m1), .pwm_clk(pwm_clk), 
            .free_m1(free_m1), .clkout_c_enable_244(clkout_c_enable_244), 
            .PWMdut_m1({PWMdut_m1}), .hallsense_m1({hallsense_m1}), .n21920(n21920), 
            .enable_m1(enable_m1), .n2798(n2798), .n2834(n2834), .n21918(n21918));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(308[13:25])
    HALL_U4 HALL_I_M2 (.clk_1mhz(clk_1mhz), .\speed_m2[0] (speed_m2[0]), 
            .hallsense_m2({hallsense_m2}), .clkout_c_enable_244(clkout_c_enable_244), 
            .clkout_c_enable_219(clkout_c_enable_219), .H_C_m2_c(H_C_m2_c), 
            .H_B_m2_c(H_B_m2_c), .H_A_m2_c(H_A_m2_c), .\speed_m2[1] (speed_m2[1]), 
            .\speed_m2[2] (speed_m2[2]), .\speed_m2[3] (speed_m2[3]), .\speed_m2[4] (speed_m2[4]), 
            .\speed_m2[5] (speed_m2[5]), .\speed_m2[6] (speed_m2[6]), .\speed_m2[7] (speed_m2[7]), 
            .\speed_m2[8] (speed_m2[8]), .\speed_m2[9] (speed_m2[9]), .\speed_m2[10] (speed_m2[10]), 
            .\speed_m2[11] (speed_m2[11]), .\speed_m2[12] (speed_m2[12]), 
            .\speed_m2[13] (speed_m2[13]), .\speed_m2[14] (speed_m2[14]), 
            .\speed_m2[15] (speed_m2[15]), .\speed_m2[16] (speed_m2[16]), 
            .\speed_m2[17] (speed_m2[17]), .\speed_m2[18] (speed_m2[18]), 
            .\speed_m2[19] (speed_m2[19]), .n22378(n22378), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(312[14:18])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    SPI SPI_I (.MISO_N_624(MISO_N_624), .clkout_c(clkout_c), .enable_m4(enable_m4), 
        .clkout_c_enable_219(clkout_c_enable_219), .speed_set_m3({speed_set_m3}), 
        .HALL_A_OUT_c_c(HALL_A_OUT_c_c), .clkout_c_enable_244(clkout_c_enable_244), 
        .HALL_B_OUT_c_c(HALL_B_OUT_c_c), .enable_m1(enable_m1), .free_m1(free_m1), 
        .hallsense_m1({hallsense_m1}), .n20053(n20053), .enable_m2(enable_m2), 
        .n21864(n21864), .enable_m3(enable_m3), .HALL_C_OUT_c_c(HALL_C_OUT_c_c), 
        .n21865(n21865), .dir_m1(dir_m1), .n2786(n2786), .n2822(n2822), 
        .hallsense_m2({hallsense_m2}), .dir_m2(dir_m2), .n2916(n2916), 
        .n2952(n2952), .speed_set_m4({speed_set_m4}), .hallsense_m3({hallsense_m3}), 
        .n21907(n21907), .dir_m3(dir_m3), .n3046(n3046), .n3082(n3082), 
        .speed_set_m2({speed_set_m2}), .n22383(n22383), .rst(rst), .\send_buffer[94] (send_buffer[94]), 
        .\send_buffer_95__N_346[94] (send_buffer_95__N_346[94]), .hallsense_m4({hallsense_m4}), 
        .dir_m4(dir_m4), .n3176(n3176), .n3212(n3212), .GND_net(GND_net), 
        .speed_set_m1({speed_set_m1}), .\speed_m1[19] (speed_m1[19]), .\speed_m2[1] (speed_m2[1]), 
        .\speed_m2[2] (speed_m2[2]), .\speed_m3[19] (speed_m3[19]), .\speed_m2[3] (speed_m2[3]), 
        .\speed_m2[0] (speed_m2[0]), .\speed_m2[4] (speed_m2[4]), .\speed_m2[5] (speed_m2[5]), 
        .\speed_m2[6] (speed_m2[6]), .\speed_m2[7] (speed_m2[7]), .\speed_m2[8] (speed_m2[8]), 
        .\speed_m2[9] (speed_m2[9]), .\speed_m2[10] (speed_m2[10]), .\speed_m2[11] (speed_m2[11]), 
        .\speed_m2[12] (speed_m2[12]), .\speed_m2[13] (speed_m2[13]), .\speed_m2[14] (speed_m2[14]), 
        .\speed_m2[15] (speed_m2[15]), .\speed_m2[16] (speed_m2[16]), .\speed_m2[17] (speed_m2[17]), 
        .\speed_m4[6] (speed_m4[6]), .\speed_m4[5] (speed_m4[5]), .\speed_m2[18] (speed_m2[18]), 
        .\speed_m2[19] (speed_m2[19]), .\speed_m1[0] (speed_m1[0]), .\speed_m1[1] (speed_m1[1]), 
        .\speed_m1[2] (speed_m1[2]), .\speed_m1[3] (speed_m1[3]), .\speed_m1[4] (speed_m1[4]), 
        .\speed_m1[5] (speed_m1[5]), .\speed_m1[6] (speed_m1[6]), .\speed_m1[7] (speed_m1[7]), 
        .\speed_m1[8] (speed_m1[8]), .\speed_m1[9] (speed_m1[9]), .\speed_m1[10] (speed_m1[10]), 
        .\speed_m1[11] (speed_m1[11]), .\speed_m1[12] (speed_m1[12]), .\speed_m1[13] (speed_m1[13]), 
        .\speed_m1[14] (speed_m1[14]), .\speed_m1[15] (speed_m1[15]), .\speed_m1[16] (speed_m1[16]), 
        .\speed_m4[8] (speed_m4[8]), .\speed_m4[7] (speed_m4[7]), .\speed_m1[17] (speed_m1[17]), 
        .\speed_m1[18] (speed_m1[18]), .\speed_m4[10] (speed_m4[10]), .\speed_m4[9] (speed_m4[9]), 
        .\speed_m4[11] (speed_m4[11]), .\speed_m4[12] (speed_m4[12]), .\speed_m4[13] (speed_m4[13]), 
        .\speed_m4[14] (speed_m4[14]), .\speed_m4[15] (speed_m4[15]), .\speed_m4[16] (speed_m4[16]), 
        .\speed_m4[17] (speed_m4[17]), .\speed_m4[18] (speed_m4[18]), .\speed_m4[19] (speed_m4[19]), 
        .\speed_m3[0] (speed_m3[0]), .\speed_m3[1] (speed_m3[1]), .\speed_m3[2] (speed_m3[2]), 
        .\speed_m3[3] (speed_m3[3]), .\speed_m3[4] (speed_m3[4]), .\speed_m3[5] (speed_m3[5]), 
        .\speed_m3[6] (speed_m3[6]), .\speed_m3[7] (speed_m3[7]), .\speed_m3[8] (speed_m3[8]), 
        .\speed_m3[9] (speed_m3[9]), .n4884(n4884), .\speed_m3[10] (speed_m3[10]), 
        .\speed_m3[11] (speed_m3[11]), .\speed_m3[12] (speed_m3[12]), .\speed_m3[13] (speed_m3[13]), 
        .\speed_m3[14] (speed_m3[14]), .\speed_m3[15] (speed_m3[15]), .\speed_m3[16] (speed_m3[16]), 
        .\speed_m3[17] (speed_m3[17]), .\speed_m3[18] (speed_m3[18]), .\speed_m4[0] (speed_m4[0]), 
        .\speed_m4[1] (speed_m4[1]), .\speed_m4[2] (speed_m4[2]), .\speed_m4[3] (speed_m4[3]), 
        .\speed_m4[4] (speed_m4[4]), .free_m4(free_m4), .n20030(n20030), 
        .free_m2(free_m2), .n20041(n20041));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(293[10:13])
    FD1P3AX start_cnt_2059__i1 (.D(n74), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i1.GSR = "DISABLED";
    HALL HALL_I_M4 (.clk_1mhz(clk_1mhz), .\speed_m4[0] (speed_m4[0]), .clkout_c_enable_244(clkout_c_enable_244), 
         .hallsense_m4({hallsense_m4}), .H_A_m4_c(H_A_m4_c), .H_B_m4_c(H_B_m4_c), 
         .H_C_m4_c(H_C_m4_c), .clkout_c_enable_219(clkout_c_enable_219), 
         .GND_net(GND_net), .\speed_m4[1] (speed_m4[1]), .\speed_m4[2] (speed_m4[2]), 
         .\speed_m4[3] (speed_m4[3]), .\speed_m4[4] (speed_m4[4]), .\speed_m4[5] (speed_m4[5]), 
         .\speed_m4[6] (speed_m4[6]), .\speed_m4[7] (speed_m4[7]), .\speed_m4[8] (speed_m4[8]), 
         .\speed_m4[9] (speed_m4[9]), .\speed_m4[10] (speed_m4[10]), .\speed_m4[11] (speed_m4[11]), 
         .\speed_m4[12] (speed_m4[12]), .\speed_m4[13] (speed_m4[13]), .\speed_m4[14] (speed_m4[14]), 
         .\speed_m4[15] (speed_m4[15]), .\speed_m4[16] (speed_m4[16]), .\speed_m4[17] (speed_m4[17]), 
         .\speed_m4[18] (speed_m4[18]), .\speed_m4[19] (speed_m4[19]), .n22378(n22378));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(332[14:18])
    \PID(16000000,160000000,10000000)  PID_I (.clk_N_683(clk_N_683), .GND_net(GND_net), 
            .n4201(n4201), .n4200(n4200), .intgOut3({Open_0, Open_1, 
            Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, 
            Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
            Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, 
            Open_21, Open_22, intgOut3[5:0]}), .backOut2({Open_23, Open_24, 
            Open_25, Open_26, Open_27, Open_28, Open_29, Open_30, 
            Open_31, Open_32, Open_33, Open_34, Open_35, Open_36, 
            Open_37, Open_38, Open_39, Open_40, Open_41, Open_42, 
            Open_43, Open_44, Open_45, backOut2[5:0]}), .backOut3({Open_46, 
            Open_47, Open_48, Open_49, Open_50, Open_51, Open_52, 
            Open_53, Open_54, Open_55, Open_56, Open_57, Open_58, 
            Open_59, Open_60, Open_61, Open_62, Open_63, Open_64, 
            Open_65, Open_66, Open_67, Open_68, backOut3[5:0]}), .\subOut_24__N_1135[0] (subOut_24__N_1135[0]), 
            .n4203(n4203), .n4202(n4202), .dir_m2(dir_m2), .dir_m3(dir_m3), 
            .dir_m1(dir_m1), .dir_m4(dir_m4), .n21851(n21851), .n21835(n21835), 
            .\speed_m4[3] (speed_m4[3]), .n4133(n4133), .\speed_m4[7] (speed_m4[7]), 
            .\speed_m4[8] (speed_m4[8]), .\speed_m4[9] (speed_m4[9]), .\speed_m4[12] (speed_m4[12]), 
            .speed_set_m2({speed_set_m2}), .speed_set_m3({speed_set_m3}), 
            .n20537(n20537), .n4204(n4204), .n10(n10), .n10_adj_1(n10_adj_1955), 
            .VCC_net(VCC_net), .n32(n32), .n10_adj_2(n10_adj_1953), .n10_adj_3(n10_adj_1950), 
            .n10_adj_4(n10_adj_1948), .n21(n21_adj_1959), .n21_adj_5(n21_adj_1957), 
            .n21_adj_6(n21_adj_1944), .n21_adj_7(n21_adj_1941), .n19454(n19454), 
            .n21_adj_8(n21), .n30(n30), .\subOut_24__N_1135[1] (subOut_24__N_1135[1]), 
            .\subOut_24__N_1135[2] (subOut_24__N_1135[2]), .\subOut_24__N_1135[3] (subOut_24__N_1135[3]), 
            .\subOut_24__N_1135[4] (subOut_24__N_1135[4]), .\subOut_24__N_1135[5] (subOut_24__N_1135[5]), 
            .\subOut_24__N_1135[6] (subOut_24__N_1135[6]), .\subOut_24__N_1135[7] (subOut_24__N_1135[7]), 
            .\subOut_24__N_1135[8] (subOut_24__N_1135[8]), .\subOut_24__N_1135[9] (subOut_24__N_1135[9]), 
            .\subOut_24__N_1135[10] (subOut_24__N_1135[10]), .\subOut_24__N_1135[11] (subOut_24__N_1135[11]), 
            .\subOut_24__N_1135[12] (subOut_24__N_1135[12]), .\subOut_24__N_1135[13] (subOut_24__N_1135[13]), 
            .\subOut_24__N_1135[14] (subOut_24__N_1135[14]), .\subOut_24__N_1135[15] (subOut_24__N_1135[15]), 
            .\subOut_24__N_1135[16] (subOut_24__N_1135[16]), .\subOut_24__N_1135[17] (subOut_24__N_1135[17]), 
            .\subOut_24__N_1135[18] (subOut_24__N_1135[18]), .\subOut_24__N_1135[19] (subOut_24__N_1135[19]), 
            .\subOut_24__N_1135[20] (subOut_24__N_1135[20]), .\subOut_24__N_1135[21] (subOut_24__N_1135[21]), 
            .\subOut_24__N_1135[24] (subOut_24__N_1135[24]), .\speed_m1[3] (speed_m1[3]), 
            .speed_set_m1({speed_set_m1}), .speed_set_m4({speed_set_m4}), 
            .\speed_m1[7] (speed_m1[7]), .\speed_m1[8] (speed_m1[8]), .\speed_m1[9] (speed_m1[9]), 
            .\speed_m1[12] (speed_m1[12]), .\speed_m1[19] (speed_m1[19]), 
            .\speed_m2[19] (speed_m2[19]), .n5(n5), .\speed_m1[1] (speed_m1[1]), 
            .\speed_m2[1] (speed_m2[1]), .\speed_m1[2] (speed_m1[2]), .\speed_m2[2] (speed_m2[2]), 
            .\speed_m1[4] (speed_m1[4]), .\speed_m2[4] (speed_m2[4]), .\speed_m1[5] (speed_m1[5]), 
            .\speed_m2[5] (speed_m2[5]), .\speed_m1[6] (speed_m1[6]), .\speed_m2[6] (speed_m2[6]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_m2[10] (speed_m2[10]), 
            .\speed_m1[11] (speed_m1[11]), .\speed_m2[11] (speed_m2[11]), 
            .\speed_m1[13] (speed_m1[13]), .\speed_m2[13] (speed_m2[13]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_m2[14] (speed_m2[14]), 
            .\speed_m1[15] (speed_m1[15]), .\speed_m2[15] (speed_m2[15]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_m2[16] (speed_m2[16]), 
            .\speed_m1[17] (speed_m1[17]), .\speed_m2[17] (speed_m2[17]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_m2[18] (speed_m2[18]), 
            .\speed_m1[0] (speed_m1[0]), .\speed_m2[0] (speed_m2[0]), .PWMdut_m4({PWMdut_m4}), 
            .PWMdut_m3({PWMdut_m3}), .\speed_m3[3] (speed_m3[3]), .\speed_m2[3] (speed_m2[3]), 
            .n20525(n20525), .\speed_m3[7] (speed_m3[7]), .\speed_m2[7] (speed_m2[7]), 
            .\speed_m3[8] (speed_m3[8]), .\speed_m2[8] (speed_m2[8]), .\speed_m3[9] (speed_m3[9]), 
            .\speed_m2[9] (speed_m2[9]), .\speed_m3[12] (speed_m3[12]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_m4[1] (speed_m4[1]), 
            .\speed_m3[1] (speed_m3[1]), .n21857(n21857), .\speed_m4[2] (speed_m4[2]), 
            .\speed_m3[2] (speed_m3[2]), .\speed_m4[4] (speed_m4[4]), .\speed_m3[4] (speed_m3[4]), 
            .\speed_m4[5] (speed_m4[5]), .\speed_m3[5] (speed_m3[5]), .\speed_m4[6] (speed_m4[6]), 
            .\speed_m3[6] (speed_m3[6]), .\speed_m4[10] (speed_m4[10]), 
            .\speed_m3[10] (speed_m3[10]), .\speed_m4[11] (speed_m4[11]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_m4[13] (speed_m4[13]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_m4[14] (speed_m4[14]), 
            .\speed_m3[14] (speed_m3[14]), .\speed_m4[15] (speed_m4[15]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_m4[16] (speed_m4[16]), 
            .\speed_m3[16] (speed_m3[16]), .\speed_m4[17] (speed_m4[17]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_m4[18] (speed_m4[18]), 
            .\speed_m3[18] (speed_m3[18]), .\speed_m4[0] (speed_m4[0]), 
            .\speed_m3[0] (speed_m3[0]), .PWMdut_m2({PWMdut_m2}), .n9(n9), 
            .PWMdut_m1({PWMdut_m1}), .n20586(n20586), .n22383(n22383), 
            .n4208(n4208), .n7(n7), .n4210(n4210), .n4209(n4209), .n4212(n4212), 
            .n4211(n4211), .n4214(n4214), .n4213(n4213), .n4216(n4216), 
            .n4215(n4215), .n4218(n4218), .n4217(n4217), .n4220(n4220), 
            .n4219(n4219), .n4222(n4222), .n4221(n4221), .n4224(n4224), 
            .n4223(n4223), .n4226(n4226), .n4225(n4225), .n4228(n4228), 
            .n4227(n4227), .n4229(n4229), .n4183(n4183), .n4182(n4182), 
            .n13(n13), .n4185(n4185), .n4184(n4184), .n13_adj_9(n13_adj_1956), 
            .n13_adj_10(n13_adj_1940), .n4187(n4187), .n4186(n4186), .n13_adj_11(n13_adj_1939), 
            .n13_adj_12(n13_adj_1943), .n4189(n4189), .n4188(n4188), .n14(n14), 
            .n4191(n4191), .n4190(n4190), .n4193(n4193), .n4192(n4192), 
            .n4195(n4195), .n4194(n4194), .n4197(n4197), .n4196(n4196), 
            .n4199(n4199), .n4198(n4198));   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(297[10:13])
    FD1P3AX start_cnt_2059__i2 (.D(n73), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i2.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i3 (.D(n72), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i3.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i4 (.D(n71), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i4.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i5 (.D(n70), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i5.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i6 (.D(n69), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i6.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i7 (.D(n68), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i7.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i8 (.D(n67), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i8.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i9 (.D(n66), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i9.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i10 (.D(n65), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i10.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i11 (.D(n64), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i11.GSR = "DISABLED";
    FD1P3AX start_cnt_2059__i12 (.D(n63), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i12.GSR = "DISABLED";
    FD1S3AX start_cnt_2059__i13 (.D(n10082), .CK(clkout_c), .Q(start_cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2059__i13.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module CLKDIV
//

module CLKDIV (clkout_c, clk_1mhz, pwm_clk, GND_net, clk_N_683);
    input clkout_c;
    output clk_1mhz;
    output pwm_clk;
    input GND_net;
    output clk_N_683;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(88[9:16])
    wire pi_clk /* synthesis is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(89[9:15])
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(30[4:14])
    
    wire mhz_buf, mhz_buf_N_68, pi_buf, pi_buf_N_69, pwm_buf, pwm_buf_N_67, 
        n12990, n12989;
    wire [4:0]count;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(41[8:13])
    
    wire n20335;
    wire [4:0]n25;
    wire [11:0]cntpi;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(42[8:13])
    wire [8:0]n41;
    
    wire n21891, n20393, n20391, n18839, n18838, n18837, n18836;
    
    FD1S3AX mhz_buf_29 (.D(mhz_buf_N_68), .CK(clkout_c), .Q(mhz_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(55[1] 79[8])
    defparam mhz_buf_29.GSR = "DISABLED";
    FD1S3AX pi_buf_30 (.D(pi_buf_N_69), .CK(clkout_c), .Q(pi_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(55[1] 79[8])
    defparam pi_buf_30.GSR = "DISABLED";
    FD1S3AX pwm_buf_32 (.D(pwm_buf_N_67), .CK(clkout_c), .Q(pwm_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(55[1] 79[8])
    defparam pwm_buf_32.GSR = "DISABLED";
    FD1S3AX clk_1mhz_33 (.D(mhz_buf), .CK(clkout_c), .Q(clk_1mhz)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(55[1] 79[8])
    defparam clk_1mhz_33.GSR = "DISABLED";
    FD1S3AX pwm_clk_34 (.D(pwm_buf), .CK(clkout_c), .Q(pwm_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(55[1] 79[8])
    defparam pwm_clk_34.GSR = "DISABLED";
    FD1S3AX pi_clk_35 (.D(pi_buf), .CK(clkout_c), .Q(pi_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(55[1] 79[8])
    defparam pi_clk_35.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(mhz_buf), .B(n12990), .Z(mhz_buf_N_68)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_200 (.A(pi_buf), .B(n12989), .Z(pi_buf_N_69)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_200.init = 16'h6666;
    LUT4 i18312_4_lut (.A(count[2]), .B(count[0]), .C(count[3]), .D(n20335), 
         .Z(n12990)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(61[5:15])
    defparam i18312_4_lut.init = 16'h0400;
    LUT4 i17510_2_lut (.A(count[4]), .B(count[1]), .Z(n20335)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17510_2_lut.init = 16'h8888;
    LUT4 i16140_1_lut (.A(count[0]), .Z(n25[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam i16140_1_lut.init = 16'h5555;
    FD1S3IX count_2060__i0 (.D(n25[0]), .CK(clkout_c), .CD(n12990), .Q(count[0]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam count_2060__i0.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i1 (.D(n41[0]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i1.GSR = "DISABLED";
    LUT4 i16163_3_lut_4_lut (.A(count[2]), .B(n21891), .C(count[3]), .D(count[4]), 
         .Z(n25[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam i16163_3_lut_4_lut.init = 16'h7f80;
    LUT4 i18309_4_lut (.A(n20393), .B(cntpi[2]), .C(n20391), .D(cntpi[7]), 
         .Z(n12989)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(66[5:16])
    defparam i18309_4_lut.init = 16'h0020;
    LUT4 i17567_3_lut (.A(cntpi[5]), .B(cntpi[3]), .C(cntpi[6]), .Z(n20393)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17567_3_lut.init = 16'h8080;
    LUT4 i17565_4_lut (.A(cntpi[1]), .B(cntpi[0]), .C(cntpi[8]), .D(cntpi[4]), 
         .Z(n20391)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17565_4_lut.init = 16'h8000;
    LUT4 pwm_buf_I_0_1_lut (.A(pwm_buf), .Z(pwm_buf_N_67)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(73[14:25])
    defparam pwm_buf_I_0_1_lut.init = 16'h5555;
    LUT4 i16145_2_lut_rep_471 (.A(count[1]), .B(count[0]), .Z(n21891)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam i16145_2_lut_rep_471.init = 16'h8888;
    LUT4 i16149_2_lut_3_lut (.A(count[1]), .B(count[0]), .C(count[2]), 
         .Z(n25[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam i16149_2_lut_3_lut.init = 16'h7878;
    LUT4 i16156_2_lut_3_lut_4_lut (.A(count[1]), .B(count[0]), .C(count[3]), 
         .D(count[2]), .Z(n25[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam i16156_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D cntpi_2061_2062_add_4_9 (.A0(cntpi[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18839), .S0(n41[7]), .S1(n41[8]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062_add_4_9.INIT0 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_9.INIT1 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_9.INJECT1_0 = "NO";
    defparam cntpi_2061_2062_add_4_9.INJECT1_1 = "NO";
    CCU2D cntpi_2061_2062_add_4_7 (.A0(cntpi[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18838), .COUT(n18839), .S0(n41[5]), .S1(n41[6]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062_add_4_7.INIT0 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_7.INIT1 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_7.INJECT1_0 = "NO";
    defparam cntpi_2061_2062_add_4_7.INJECT1_1 = "NO";
    CCU2D cntpi_2061_2062_add_4_5 (.A0(cntpi[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18837), .COUT(n18838), .S0(n41[3]), .S1(n41[4]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062_add_4_5.INIT0 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_5.INIT1 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_5.INJECT1_0 = "NO";
    defparam cntpi_2061_2062_add_4_5.INJECT1_1 = "NO";
    CCU2D cntpi_2061_2062_add_4_3 (.A0(cntpi[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18836), .COUT(n18837), .S0(n41[1]), .S1(n41[2]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062_add_4_3.INIT0 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_3.INIT1 = 16'hfaaa;
    defparam cntpi_2061_2062_add_4_3.INJECT1_0 = "NO";
    defparam cntpi_2061_2062_add_4_3.INJECT1_1 = "NO";
    CCU2D cntpi_2061_2062_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18836), .S1(n41[0]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062_add_4_1.INIT0 = 16'hF000;
    defparam cntpi_2061_2062_add_4_1.INIT1 = 16'h0555;
    defparam cntpi_2061_2062_add_4_1.INJECT1_0 = "NO";
    defparam cntpi_2061_2062_add_4_1.INJECT1_1 = "NO";
    LUT4 i16142_2_lut (.A(count[1]), .B(count[0]), .Z(n25[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam i16142_2_lut.init = 16'h6666;
    INV i18552 (.A(pi_clk), .Z(clk_N_683));
    FD1S3IX cntpi_2061_2062__i2 (.D(n41[1]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i2.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i3 (.D(n41[2]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i3.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i4 (.D(n41[3]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i4.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i5 (.D(n41[4]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i5.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i6 (.D(n41[5]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i6.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i7 (.D(n41[6]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i7.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i8 (.D(n41[7]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i8.GSR = "DISABLED";
    FD1S3IX cntpi_2061_2062__i9 (.D(n41[8]), .CK(clkout_c), .CD(n12989), 
            .Q(cntpi[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(57[11:16])
    defparam cntpi_2061_2062__i9.GSR = "DISABLED";
    FD1S3IX count_2060__i1 (.D(n25[1]), .CK(clkout_c), .CD(n12990), .Q(count[1]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam count_2060__i1.GSR = "DISABLED";
    FD1S3IX count_2060__i2 (.D(n25[2]), .CK(clkout_c), .CD(n12990), .Q(count[2]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam count_2060__i2.GSR = "DISABLED";
    FD1S3IX count_2060__i3 (.D(n25[3]), .CK(clkout_c), .CD(n12990), .Q(count[3]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam count_2060__i3.GSR = "DISABLED";
    FD1S3IX count_2060__i4 (.D(n25[4]), .CK(clkout_c), .CD(n12990), .Q(count[4]));   // c:/users/gebruiker/workspace/lattice/final code software/clockdivider.vhd(56[11:16])
    defparam count_2060__i4.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION_U8
//

module COMMUTATION_U8 (MB_m1_c_0, clkout_c, MC_m1_c_0, MA_m1_c_0, LED1_c, 
            MA_m1_c_1, n20053, n2880, MC_m1_c_1, n2834, n2822, MB_m1_c_1, 
            n2798, n2786, enable_m1, n21920, PWM_m1, n21918, n21917, 
            free_m1);
    output MB_m1_c_0;
    input clkout_c;
    output MC_m1_c_0;
    output MA_m1_c_0;
    output LED1_c;
    output MA_m1_c_1;
    input n20053;
    input n2880;
    output MC_m1_c_1;
    input n2834;
    input n2822;
    output MB_m1_c_1;
    input n2798;
    input n2786;
    input enable_m1;
    input n21920;
    input PWM_m1;
    input n21918;
    input n21917;
    input free_m1;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n19076, n19075, n20054, clkout_c_enable_4;
    
    FD1S3IX MospairB_i1 (.D(n19076), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n19075), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n20054), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_4), .CK(clkout_c), 
            .Q(LED1_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    FD1S3IX MospairA_i2 (.D(n2880), .CK(clkout_c), .CD(n20053), .Q(MA_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n2822), .CK(clkout_c), .CD(n2834), .Q(MC_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2786), .CK(clkout_c), .CD(n2798), .Q(MB_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i10310_1_lut (.A(enable_m1), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i10310_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2786), .B(n21920), .C(PWM_m1), .Z(n19076)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_199 (.A(n2822), .B(n21918), .C(PWM_m1), .Z(n19075)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_199.init = 16'hbfbf;
    LUT4 i18325_3_lut (.A(n20053), .B(PWM_m1), .C(n21917), .Z(n20054)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i18325_3_lut.init = 16'hbfbf;
    LUT4 i18388_2_lut (.A(free_m1), .B(enable_m1), .Z(clkout_c_enable_4)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i18388_2_lut.init = 16'h7777;
    
endmodule
//
// Verilog Description of module COMMUTATION_U7
//

module COMMUTATION_U7 (MB_m2_c_0, clkout_c, MC_m2_c_0, MA_m2_c_0, LED2_c, 
            MA_m2_c_1, n20041, n3010, MC_m2_c_1, n2964, n2952, MB_m2_c_1, 
            n2928, n2916, enable_m2, n21913, PWM_m2, n21911, n21910, 
            free_m2);
    output MB_m2_c_0;
    input clkout_c;
    output MC_m2_c_0;
    output MA_m2_c_0;
    output LED2_c;
    output MA_m2_c_1;
    input n20041;
    input n3010;
    output MC_m2_c_1;
    input n2964;
    input n2952;
    output MB_m2_c_1;
    input n2928;
    input n2916;
    input enable_m2;
    input n21913;
    input PWM_m2;
    input n21911;
    input n21910;
    input free_m2;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n19074, n19073, n20042, clkout_c_enable_5;
    
    FD1S3IX MospairB_i1 (.D(n19074), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n19073), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n20042), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_5), .CK(clkout_c), 
            .Q(LED2_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    FD1S3IX MospairA_i2 (.D(n3010), .CK(clkout_c), .CD(n20041), .Q(MA_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n2952), .CK(clkout_c), .CD(n2964), .Q(MC_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2916), .CK(clkout_c), .CD(n2928), .Q(MB_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i10311_1_lut (.A(enable_m2), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i10311_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2916), .B(n21913), .C(PWM_m2), .Z(n19074)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_198 (.A(n2952), .B(n21911), .C(PWM_m2), .Z(n19073)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_198.init = 16'hbfbf;
    LUT4 i18322_3_lut (.A(n20041), .B(PWM_m2), .C(n21910), .Z(n20042)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i18322_3_lut.init = 16'hbfbf;
    LUT4 i18385_2_lut (.A(free_m2), .B(enable_m2), .Z(clkout_c_enable_5)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i18385_2_lut.init = 16'h7777;
    
endmodule
//
// Verilog Description of module COMMUTATION_U6
//

module COMMUTATION_U6 (MB_m3_c_0, clkout_c, MC_m3_c_0, MA_m3_c_0, LED3_c, 
            MA_m3_c_1, n20051, n3140, MC_m3_c_1, n3094, n3082, MB_m3_c_1, 
            n3058, n3046, enable_m3, n21908, PWM_m3, n21906, n21905, 
            free_m3);
    output MB_m3_c_0;
    input clkout_c;
    output MC_m3_c_0;
    output MA_m3_c_0;
    output LED3_c;
    output MA_m3_c_1;
    input n20051;
    input n3140;
    output MC_m3_c_1;
    input n3094;
    input n3082;
    output MB_m3_c_1;
    input n3058;
    input n3046;
    input enable_m3;
    input n21908;
    input PWM_m3;
    input n21906;
    input n21905;
    input free_m3;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n19072, n19063, n20052, clkout_c_enable_8;
    
    FD1S3IX MospairB_i1 (.D(n19072), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n19063), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n20052), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_8), .CK(clkout_c), 
            .Q(LED3_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    FD1S3IX MospairA_i2 (.D(n3140), .CK(clkout_c), .CD(n20051), .Q(MA_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3082), .CK(clkout_c), .CD(n3094), .Q(MC_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3046), .CK(clkout_c), .CD(n3058), .Q(MB_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i10312_1_lut (.A(enable_m3), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i10312_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3046), .B(n21908), .C(PWM_m3), .Z(n19072)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_197 (.A(n3082), .B(n21906), .C(PWM_m3), .Z(n19063)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_197.init = 16'hbfbf;
    LUT4 i18264_3_lut (.A(n20051), .B(PWM_m3), .C(n21905), .Z(n20052)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i18264_3_lut.init = 16'hbfbf;
    LUT4 i18382_2_lut (.A(free_m3), .B(enable_m3), .Z(clkout_c_enable_8)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i18382_2_lut.init = 16'h7777;
    
endmodule
//
// Verilog Description of module COMMUTATION
//

module COMMUTATION (MB_m4_c_0, clkout_c, MC_m4_c_0, MA_m4_c_0, LED4_c, 
            MA_m4_c_1, n20030, n3270, MC_m4_c_1, n3224, n3212, MB_m4_c_1, 
            n3188, n3176, enable_m4, n21902, PWM_m4, n21900, n21899, 
            free_m4);
    output MB_m4_c_0;
    input clkout_c;
    output MC_m4_c_0;
    output MA_m4_c_0;
    output LED4_c;
    output MA_m4_c_1;
    input n20030;
    input n3270;
    output MC_m4_c_1;
    input n3224;
    input n3212;
    output MB_m4_c_1;
    input n3188;
    input n3176;
    input enable_m4;
    input n21902;
    input PWM_m4;
    input n21900;
    input n21899;
    input free_m4;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n19137, n19136, n20031, clkout_c_enable_10;
    
    FD1S3IX MospairB_i1 (.D(n19137), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n19136), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n20031), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_10), .CK(clkout_c), 
            .Q(LED4_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    FD1S3IX MospairA_i2 (.D(n3270), .CK(clkout_c), .CD(n20030), .Q(MA_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3212), .CK(clkout_c), .CD(n3224), .Q(MC_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3176), .CK(clkout_c), .CD(n3188), .Q(MB_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i10316_1_lut (.A(enable_m4), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i10316_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3176), .B(n21902), .C(PWM_m4), .Z(n19137)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_196 (.A(n3212), .B(n21900), .C(PWM_m4), .Z(n19136)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_196.init = 16'hbfbf;
    LUT4 i18400_3_lut (.A(n20030), .B(PWM_m4), .C(n21899), .Z(n20031)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i18400_3_lut.init = 16'hbfbf;
    LUT4 i18379_2_lut (.A(free_m4), .B(enable_m4), .Z(clkout_c_enable_10)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i18379_2_lut.init = 16'h7777;
    
endmodule
//
// Verilog Description of module HALL_U3
//

module HALL_U3 (clk_1mhz, \speed_m3[0] , hallsense_m3, clkout_c_enable_244, 
            H_A_m3_c, H_B_m3_c, H_C_m3_c, clkout_c_enable_219, \speed_m3[1] , 
            \speed_m3[2] , \speed_m3[3] , \speed_m3[4] , \speed_m3[5] , 
            \speed_m3[6] , \speed_m3[7] , \speed_m3[8] , \speed_m3[9] , 
            \speed_m3[10] , \speed_m3[11] , \speed_m3[12] , \speed_m3[13] , 
            \speed_m3[14] , \speed_m3[15] , \speed_m3[16] , \speed_m3[17] , 
            \speed_m3[18] , \speed_m3[19] , n22378, GND_net);
    input clk_1mhz;
    output \speed_m3[0] ;
    output [2:0]hallsense_m3;
    input clkout_c_enable_244;
    input H_A_m3_c;
    input H_B_m3_c;
    input H_C_m3_c;
    input clkout_c_enable_219;
    output \speed_m3[1] ;
    output \speed_m3[2] ;
    output \speed_m3[3] ;
    output \speed_m3[4] ;
    output \speed_m3[5] ;
    output \speed_m3[6] ;
    output \speed_m3[7] ;
    output \speed_m3[8] ;
    output \speed_m3[9] ;
    output \speed_m3[10] ;
    output \speed_m3[11] ;
    output \speed_m3[12] ;
    output \speed_m3[13] ;
    output \speed_m3[14] ;
    output \speed_m3[15] ;
    output \speed_m3[16] ;
    output \speed_m3[17] ;
    output \speed_m3[18] ;
    output \speed_m3[19] ;
    input n22378;
    input GND_net;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(62[10:22])
    
    wire stable_counting, n33;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_lat, hall1_lat, hall2_lat, hall3_old, hall1_old, hall2_old;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_102, n4332;
    wire [19:0]n7;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(60[10:15])
    
    wire n12, n20043, n21841, n21855;
    wire [6:0]n83;
    
    wire n20134, n20139, n20136, n20135, n20138, n20137, stable_counting_N_1758, 
        n21874, n21875, stable_counting_N_1746, n20_adj_1935, n21828, 
        n20309, n12980;
    wire [6:0]stable_counting_N_1759;
    
    wire n21854, n20243, n16208, n20_adj_1936, n16_adj_1937, n18_adj_1938, 
        n20369, n4, n21856, n21909, n21842, n18743, n18742, n18741, 
        n18740, n18739, n18738, n18737, n18736, n18735, n18734, 
        n20097, n20094, n6, n20399;
    
    FD1P3AX stable_count__i0 (.D(n33), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m3_c), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m3_c), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m3_c), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3IX speedt__i0 (.D(n7[0]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    LUT4 i6_4_lut_rep_421 (.A(count[13]), .B(n12), .C(count[7]), .D(n20043), 
         .Z(n21841)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i6_4_lut_rep_421.init = 16'hfeff;
    LUT4 i2447_3_lut_4_lut (.A(stable_count[4]), .B(n21855), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n83[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2447_3_lut_4_lut.init = 16'h7f80;
    FD1P3AX stable_count__i6 (.D(n20134), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3AX stable_count__i5 (.D(n20139), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3AX stable_count__i4 (.D(n20136), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3AX stable_count__i3 (.D(n20135), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3AX stable_count__i2 (.D(n20138), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3AX stable_count__i1 (.D(n20137), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    LUT4 mux_28_i2_4_lut (.A(n7[1]), .B(speedt[1]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hac0a;
    LUT4 mux_28_i3_4_lut (.A(n7[2]), .B(speedt[2]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hac0a;
    LUT4 mux_28_i4_4_lut (.A(n7[3]), .B(speedt[3]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hac0a;
    LUT4 mux_28_i5_4_lut (.A(n7[4]), .B(speedt[4]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hac0a;
    LUT4 mux_28_i6_4_lut (.A(n7[5]), .B(speedt[5]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hac0a;
    LUT4 mux_28_i7_4_lut (.A(n7[6]), .B(speedt[6]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hac0a;
    LUT4 mux_28_i8_4_lut (.A(n7[7]), .B(speedt[7]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hac0a;
    LUT4 mux_28_i9_4_lut (.A(n7[8]), .B(speedt[8]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hac0a;
    LUT4 mux_28_i10_4_lut (.A(n7[9]), .B(speedt[9]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hac0a;
    LUT4 mux_28_i11_4_lut (.A(n7[10]), .B(speedt[10]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hac0a;
    LUT4 mux_28_i12_4_lut (.A(n7[11]), .B(speedt[11]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hac0a;
    LUT4 mux_28_i13_4_lut (.A(n7[12]), .B(speedt[12]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hac0a;
    LUT4 mux_28_i14_4_lut (.A(n7[13]), .B(speedt[13]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hac0a;
    LUT4 mux_28_i15_4_lut (.A(n7[14]), .B(speedt[14]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hac0a;
    LUT4 mux_28_i16_4_lut (.A(n7[15]), .B(speedt[15]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hac0a;
    LUT4 mux_28_i17_4_lut (.A(n7[16]), .B(speedt[16]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hac0a;
    LUT4 mux_28_i18_4_lut (.A(n7[17]), .B(speedt[17]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hac0a;
    LUT4 mux_28_i19_4_lut (.A(n7[18]), .B(speedt[18]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hac0a;
    LUT4 mux_28_i20_4_lut (.A(n7[19]), .B(speedt[19]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hac0a;
    LUT4 i1_3_lut_4_lut (.A(stable_count[3]), .B(n21874), .C(n21875), 
         .D(stable_counting_N_1746), .Z(n20_adj_1935)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (B (D)+!B ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i1_3_lut_4_lut.init = 16'hff09;
    LUT4 i2440_2_lut_rep_408_3_lut_4_lut (.A(stable_count[3]), .B(n21874), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21828)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2440_2_lut_rep_408_3_lut_4_lut.init = 16'h78f0;
    LUT4 i17485_2_lut_3_lut_4_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21874), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n20309)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i17485_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h7ff8;
    LUT4 i18391_2_lut_3_lut_3_lut_4_lut (.A(stable_count[0]), .B(stable_counting_N_1746), 
         .C(stable_counting), .D(stable_counting_N_1758), .Z(n33)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;
    defparam i18391_2_lut_3_lut_3_lut_4_lut.init = 16'h0111;
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n7[1]), .CK(clk_1mhz), .CD(n12980), .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n7[2]), .CK(clk_1mhz), .CD(n12980), .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n7[3]), .CK(clk_1mhz), .CD(n12980), .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n7[4]), .CK(clk_1mhz), .CD(n12980), .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n7[5]), .CK(clk_1mhz), .CD(n12980), .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n7[6]), .CK(clk_1mhz), .CD(n12980), .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n7[7]), .CK(clk_1mhz), .CD(n12980), .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n7[8]), .CK(clk_1mhz), .CD(n12980), .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n7[9]), .CK(clk_1mhz), .CD(n12980), .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n7[10]), .CK(clk_1mhz), .CD(n12980), .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n7[11]), .CK(clk_1mhz), .CD(n12980), .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n7[12]), .CK(clk_1mhz), .CD(n12980), .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n7[13]), .CK(clk_1mhz), .CD(n12980), .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n7[14]), .CK(clk_1mhz), .CD(n12980), .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n7[15]), .CK(clk_1mhz), .CD(n12980), .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n7[16]), .CK(clk_1mhz), .CD(n12980), .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n7[17]), .CK(clk_1mhz), .CD(n12980), .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n7[18]), .CK(clk_1mhz), .CD(n12980), .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n7[19]), .CK(clk_1mhz), .CD(n12980), .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(stable_counting_N_1759[1]), .B(n21854), .C(n20309), 
         .D(n20243), .Z(stable_counting_N_1758)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[7:23])
    defparam i3_4_lut.init = 16'h0002;
    LUT4 i15_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n83[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(62[10:22])
    defparam i15_2_lut.init = 16'h6666;
    LUT4 mux_28_i1_4_lut (.A(n7[0]), .B(speedt[0]), .C(stable_counting_N_1758), 
         .D(n21841), .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hac0a;
    LUT4 i5_4_lut (.A(count[6]), .B(n16208), .C(count[15]), .D(count[11]), 
         .Z(n12)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_188 (.A(count[12]), .B(count[10]), .C(count[0]), 
         .D(count[8]), .Z(n16208)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i3_4_lut_adj_188.init = 16'hfffe;
    LUT4 i10_4_lut (.A(count[14]), .B(n20_adj_1936), .C(n16_adj_1937), 
         .D(count[1]), .Z(n20043)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i10_4_lut.init = 16'h8000;
    LUT4 i9_4_lut (.A(count[2]), .B(n18_adj_1938), .C(count[16]), .D(count[19]), 
         .Z(n20_adj_1936)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i5_2_lut (.A(count[4]), .B(count[3]), .Z(n16_adj_1937)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i5_2_lut.init = 16'h8888;
    LUT4 i7_4_lut (.A(count[18]), .B(count[9]), .C(count[5]), .D(count[17]), 
         .Z(n18_adj_1938)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i7_4_lut.init = 16'h8000;
    FD1S3IX count__i0 (.D(n7[0]), .CK(clk_1mhz), .CD(n12980), .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22378), .SP(stable_counting_N_1746), 
            .CD(n20369), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3IX speedt__i1 (.D(n7[1]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(hall2_old), .B(hall1_old), .C(hall2_lat), .D(hall1_lat), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(92[7:87])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i17543_3_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(stable_counting_N_1758), .Z(n20369)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i17543_3_lut.init = 16'hc8c8;
    FD1P3IX speedt__i2 (.D(n7[2]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n7[3]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n7[4]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n7[5]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n7[6]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n7[7]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n7[8]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n7[9]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n7[10]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n7[11]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n7[12]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n7[13]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n7[14]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n7[15]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n7[16]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n7[17]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n7[18]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n7[19]), .SP(clk_1mhz_enable_102), .CD(n4332), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_453 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_453.init = 16'hdede;
    LUT4 i13432_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .D(n83[1]), 
         .Z(stable_counting_N_1759[1])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i13432_2_lut_4_lut.init = 16'h2100;
    LUT4 i1_2_lut_rep_436_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), 
         .D(stable_count[0]), .Z(n21856)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_436_4_lut.init = 16'hffde;
    LUT4 i2433_2_lut_rep_422_3_lut_4_lut (.A(stable_count[2]), .B(n21909), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21842)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2433_2_lut_rep_422_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18743), 
          .S0(n7[19]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18742), .COUT(n18743), .S0(n7[17]), .S1(n7[18]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18741), .COUT(n18742), .S0(n7[15]), .S1(n7[16]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18740), .COUT(n18741), .S0(n7[13]), .S1(n7[14]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18739), .COUT(n18740), .S0(n7[11]), .S1(n7[12]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18738), .COUT(n18739), .S0(n7[9]), .S1(n7[10]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18737), 
          .COUT(n18738), .S0(n7[7]), .S1(n7[8]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18736), 
          .COUT(n18737), .S0(n7[5]), .S1(n7[6]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18735), 
          .COUT(n18736), .S0(n7[3]), .S1(n7[4]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18734), 
          .COUT(n18735), .S0(n7[1]), .S1(n7[2]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18734), 
          .S1(n7[0]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21841), .Z(clk_1mhz_enable_102)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n83[1]), .D(stable_counting_N_1746), .Z(n20137)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_189 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n83[6]), .D(stable_counting_N_1746), .Z(n20134)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_189.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_190 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21828), .D(stable_counting_N_1746), .Z(n20139)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_190.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_191 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21854), .D(stable_counting_N_1746), .Z(n20135)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_191.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_192 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21842), .D(stable_counting_N_1746), .Z(n20136)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_192.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_193 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21875), .D(stable_counting_N_1746), .Z(n20138)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_193.init = 16'h0070;
    LUT4 i1_2_lut_rep_489 (.A(stable_count[0]), .B(stable_count[1]), .Z(n21909)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_rep_489.init = 16'h8888;
    LUT4 i2421_2_lut_rep_454_3_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[2]), .Z(n21874)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i2421_2_lut_rep_454_3_lut.init = 16'h8080;
    LUT4 i2426_2_lut_rep_434_3_lut_4_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21854)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i2426_2_lut_rep_434_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2428_2_lut_rep_435_3_lut_4_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21855)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i2428_2_lut_rep_435_3_lut_4_lut.init = 16'h8000;
    LUT4 i2419_2_lut_rep_455_3_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[2]), .Z(n21875)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i2419_2_lut_rep_455_3_lut.init = 16'h7878;
    LUT4 i17419_3_lut_4_lut_4_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(n83[6]), .D(stable_count[2]), .Z(n20243)) /* synthesis lut_function=((B (C+!(D))+!B (C+(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i17419_3_lut_4_lut_4_lut.init = 16'hf7fd;
    LUT4 i2_3_lut (.A(n20097), .B(stable_counting), .C(n20043), .Z(n4332)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i4_4_lut (.A(count[7]), .B(n20094), .C(stable_counting_N_1759[1]), 
         .D(n6), .Z(n20097)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i4_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_194 (.A(n21856), .B(count[13]), .C(n20399), .D(n20_adj_1935), 
         .Z(n20094)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_4_lut_adj_194.init = 16'h0200;
    LUT4 i1_4_lut_adj_195 (.A(n16208), .B(n83[6]), .C(stable_counting_N_1746), 
         .D(n20309), .Z(n6)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+!(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_4_lut_adj_195.init = 16'h5051;
    LUT4 i17573_4_lut (.A(n12980), .B(count[15]), .C(count[6]), .D(count[11]), 
         .Z(n20399)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i17573_4_lut.init = 16'hfffd;
    LUT4 i18274_2_lut_3_lut_3_lut (.A(n21841), .B(stable_counting_N_1758), 
         .C(stable_counting), .Z(n12980)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i18274_2_lut_3_lut_3_lut.init = 16'hd5d5;
    
endmodule
//
// Verilog Description of module PWMGENERATOR
//

module PWMGENERATOR (PWM_m4, pwm_clk, free_m4, clkout_c_enable_244, 
            PWMdut_m4, GND_net, hallsense_m4, n21900, enable_m4, n3224, 
            n21902, n3188);
    output PWM_m4;
    input pwm_clk;
    output free_m4;
    input clkout_c_enable_244;
    input [9:0]PWMdut_m4;
    input GND_net;
    input [2:0]hallsense_m4;
    output n21900;
    input enable_m4;
    output n3224;
    output n21902;
    output n3188;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_1805, free_N_1817, n10, n7, n10_adj_1932, n10960, 
        n9;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(41[10:13])
    
    wire n12985;
    wire [9:0]n45;
    
    wire n20409, n6, n20383, n18805, n18804, n18803, n18802, n18801, 
        n3688, n18785, n14, n10_adj_1933, n18784, n18783, n18782, 
        n18781;
    
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m4)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=338, LSE_RLINE=338 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_244), .CK(pwm_clk), 
            .Q(free_m4));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(PWMdut_m4[5]), .B(PWMdut_m4[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_1932), .B(PWMdut_m4[9]), .C(PWMdut_m4[8]), 
         .D(PWMdut_m4[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2257_3_lut (.A(n10960), .B(PWMdut_m4[4]), .C(PWMdut_m4[3]), 
         .Z(n10_adj_1932)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2257_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    FD1S3IX cnt_2068__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12985), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i0.GSR = "ENABLED";
    LUT4 i18297_4_lut (.A(cnt[2]), .B(n20409), .C(cnt[1]), .D(n6), .Z(n12985)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(73[6:16])
    defparam i18297_4_lut.init = 16'h0004;
    LUT4 i17583_3_lut (.A(cnt[6]), .B(n20383), .C(cnt[8]), .Z(n20409)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17583_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[4]), .B(cnt[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i17557_4_lut (.A(cnt[7]), .B(cnt[5]), .C(cnt[9]), .D(cnt[3]), 
         .Z(n20383)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17557_4_lut.init = 16'h8000;
    CCU2D cnt_2068_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18805), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2068_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2068_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2068_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2068_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18804), 
          .COUT(n18805), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2068_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2068_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2068_add_4_9.INJECT1_1 = "NO";
    FD1S3IX cnt_2068__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12985), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i1.GSR = "ENABLED";
    CCU2D cnt_2068_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18803), 
          .COUT(n18804), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2068_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2068_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2068_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2068_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18802), 
          .COUT(n18803), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2068_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2068_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2068_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2068_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18801), 
          .COUT(n18802), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2068_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2068_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2068_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2068_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18801), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2068_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2068_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2068_add_4_1.INJECT1_1 = "NO";
    LUT4 i1798_1_lut (.A(n3688), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1798_1_lut.init = 16'h5555;
    CCU2D sub_1796_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m4[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18785), .S1(n3688));
    defparam sub_1796_add_2_11.INIT0 = 16'h5999;
    defparam sub_1796_add_2_11.INIT1 = 16'h0000;
    defparam sub_1796_add_2_11.INJECT1_0 = "NO";
    defparam sub_1796_add_2_11.INJECT1_1 = "NO";
    LUT4 i18294_4_lut (.A(PWMdut_m4[5]), .B(n14), .C(n10_adj_1933), .D(PWMdut_m4[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i18294_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m4[9]), .B(PWMdut_m4[3]), .C(PWMdut_m4[4]), 
         .D(n10960), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[7]), .Z(n10_adj_1933)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    CCU2D sub_1796_add_2_9 (.A0(PWMdut_m4[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m4[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18784), 
          .COUT(n18785));
    defparam sub_1796_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1796_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1796_add_2_9.INJECT1_0 = "NO";
    defparam sub_1796_add_2_9.INJECT1_1 = "NO";
    LUT4 i2_3_lut_adj_187 (.A(PWMdut_m4[2]), .B(PWMdut_m4[1]), .C(PWMdut_m4[0]), 
         .Z(n10960)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_187.init = 16'hfefe;
    CCU2D sub_1796_add_2_7 (.A0(PWMdut_m4[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m4[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18783), 
          .COUT(n18784));
    defparam sub_1796_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1796_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1796_add_2_7.INJECT1_0 = "NO";
    defparam sub_1796_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_5 (.A0(PWMdut_m4[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m4[4]), .C1(n9), .D1(n10), .CIN(n18782), 
          .COUT(n18783));
    defparam sub_1796_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1796_add_2_5.INIT1 = 16'h5999;
    defparam sub_1796_add_2_5.INJECT1_0 = "NO";
    defparam sub_1796_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m4[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m4[2]), .C1(n9), .D1(n10), .CIN(n18781), 
          .COUT(n18782));
    defparam sub_1796_add_2_3.INIT0 = 16'h5999;
    defparam sub_1796_add_2_3.INIT1 = 16'h5999;
    defparam sub_1796_add_2_3.INJECT1_0 = "NO";
    defparam sub_1796_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m4[0]), .C1(n9), .D1(n10), 
          .COUT(n18781));
    defparam sub_1796_add_2_1.INIT0 = 16'h0000;
    defparam sub_1796_add_2_1.INIT1 = 16'h5999;
    defparam sub_1796_add_2_1.INJECT1_0 = "NO";
    defparam sub_1796_add_2_1.INJECT1_1 = "NO";
    LUT4 i1722_3_lut_rep_480 (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .Z(n21900)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1722_3_lut_rep_480.init = 16'h1414;
    LUT4 i18367_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .D(enable_m4), .Z(n3224)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18367_2_lut_4_lut.init = 16'hebff;
    LUT4 i1692_3_lut_rep_482 (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .Z(n21902)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1692_3_lut_rep_482.init = 16'h1414;
    LUT4 i18364_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .D(enable_m4), .Z(n3188)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18364_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2068__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12985), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i2.GSR = "ENABLED";
    FD1S3IX cnt_2068__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12985), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i3.GSR = "ENABLED";
    FD1S3IX cnt_2068__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12985), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i4.GSR = "ENABLED";
    FD1S3IX cnt_2068__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12985), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i5.GSR = "ENABLED";
    FD1S3IX cnt_2068__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12985), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i6.GSR = "ENABLED";
    FD1S3IX cnt_2068__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12985), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i7.GSR = "ENABLED";
    FD1S3IX cnt_2068__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12985), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i8.GSR = "ENABLED";
    FD1S3IX cnt_2068__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12985), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2068__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U0
//

module PWMGENERATOR_U0 (PWM_m3, pwm_clk, free_m3, clkout_c_enable_219, 
            PWMdut_m3, GND_net, hallsense_m3, n21906, enable_m3, n3094, 
            n21907, n20051, n21908, n3058);
    output PWM_m3;
    input pwm_clk;
    output free_m3;
    input clkout_c_enable_219;
    input [9:0]PWMdut_m3;
    input GND_net;
    input [2:0]hallsense_m3;
    output n21906;
    input enable_m3;
    output n3094;
    output n21907;
    output n20051;
    output n21908;
    output n3058;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_1805, free_N_1817, n10, n7, n10_adj_1930, n10962, 
        n9, n18810;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(41[10:13])
    wire [9:0]n45;
    
    wire n18809, n18808, n18807, n18806, n12986, n20401, n6, n20355, 
        n3675, n18790, n18789, n18788, n18787, n18786, n14, n10_adj_1931;
    
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m3)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=328, LSE_RLINE=328 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_219), .CK(pwm_clk), 
            .Q(free_m3));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(PWMdut_m3[5]), .B(PWMdut_m3[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_1930), .B(PWMdut_m3[9]), .C(PWMdut_m3[8]), 
         .D(PWMdut_m3[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2260_3_lut (.A(n10962), .B(PWMdut_m3[4]), .C(PWMdut_m3[3]), 
         .Z(n10_adj_1930)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2260_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D cnt_2067_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18810), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2067_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18809), 
          .COUT(n18810), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18808), 
          .COUT(n18809), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18807), 
          .COUT(n18808), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18806), 
          .COUT(n18807), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_3.INJECT1_1 = "NO";
    FD1S3IX cnt_2067__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12986), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i0.GSR = "ENABLED";
    LUT4 i18300_4_lut (.A(cnt[0]), .B(n20401), .C(cnt[2]), .D(n6), .Z(n12986)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(73[6:16])
    defparam i18300_4_lut.init = 16'h0004;
    LUT4 i17575_3_lut (.A(cnt[7]), .B(n20355), .C(cnt[3]), .Z(n20401)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17575_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i17530_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n20355)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17530_4_lut.init = 16'h8000;
    CCU2D cnt_2067_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18806), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2067_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2067_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_1.INJECT1_1 = "NO";
    LUT4 i1796_1_lut (.A(n3675), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1796_1_lut.init = 16'h5555;
    CCU2D sub_1794_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m3[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18790), .S1(n3675));
    defparam sub_1794_add_2_11.INIT0 = 16'h5999;
    defparam sub_1794_add_2_11.INIT1 = 16'h0000;
    defparam sub_1794_add_2_11.INJECT1_0 = "NO";
    defparam sub_1794_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_9 (.A0(PWMdut_m3[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m3[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18789), 
          .COUT(n18790));
    defparam sub_1794_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1794_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1794_add_2_9.INJECT1_0 = "NO";
    defparam sub_1794_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_7 (.A0(PWMdut_m3[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m3[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18788), 
          .COUT(n18789));
    defparam sub_1794_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1794_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1794_add_2_7.INJECT1_0 = "NO";
    defparam sub_1794_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_5 (.A0(PWMdut_m3[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m3[4]), .C1(n9), .D1(n10), .CIN(n18787), 
          .COUT(n18788));
    defparam sub_1794_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1794_add_2_5.INIT1 = 16'h5999;
    defparam sub_1794_add_2_5.INJECT1_0 = "NO";
    defparam sub_1794_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m3[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m3[2]), .C1(n9), .D1(n10), .CIN(n18786), 
          .COUT(n18787));
    defparam sub_1794_add_2_3.INIT0 = 16'h5999;
    defparam sub_1794_add_2_3.INIT1 = 16'h5999;
    defparam sub_1794_add_2_3.INJECT1_0 = "NO";
    defparam sub_1794_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m3[0]), .C1(n9), .D1(n10), 
          .COUT(n18786));
    defparam sub_1794_add_2_1.INIT0 = 16'h0000;
    defparam sub_1794_add_2_1.INIT1 = 16'h5999;
    defparam sub_1794_add_2_1.INJECT1_0 = "NO";
    defparam sub_1794_add_2_1.INJECT1_1 = "NO";
    LUT4 i18279_4_lut (.A(PWMdut_m3[5]), .B(n14), .C(n10_adj_1931), .D(PWMdut_m3[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i18279_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m3[9]), .B(PWMdut_m3[3]), .C(PWMdut_m3[4]), 
         .D(n10962), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[7]), .Z(n10_adj_1931)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_186 (.A(PWMdut_m3[2]), .B(PWMdut_m3[1]), .C(PWMdut_m3[0]), 
         .Z(n10962)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_186.init = 16'hfefe;
    LUT4 i1630_3_lut_rep_486 (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .Z(n21906)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1630_3_lut_rep_486.init = 16'h1414;
    LUT4 i18357_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .D(enable_m3), .Z(n3094)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18357_2_lut_4_lut.init = 16'hebff;
    LUT4 i1_2_lut_rep_487 (.A(enable_m3), .B(free_m3), .Z(n21907)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1_2_lut_rep_487.init = 16'h2222;
    LUT4 i18361_3_lut_4_lut (.A(enable_m3), .B(free_m3), .C(hallsense_m3[2]), 
         .D(hallsense_m3[0]), .Z(n20051)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18361_3_lut_4_lut.init = 16'hfddf;
    LUT4 i1600_3_lut_rep_488 (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .Z(n21908)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1600_3_lut_rep_488.init = 16'h1414;
    LUT4 i18354_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .D(enable_m3), .Z(n3058)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18354_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2067__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12986), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i1.GSR = "ENABLED";
    FD1S3IX cnt_2067__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12986), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i2.GSR = "ENABLED";
    FD1S3IX cnt_2067__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12986), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i3.GSR = "ENABLED";
    FD1S3IX cnt_2067__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12986), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i4.GSR = "ENABLED";
    FD1S3IX cnt_2067__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12986), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i5.GSR = "ENABLED";
    FD1S3IX cnt_2067__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12986), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i6.GSR = "ENABLED";
    FD1S3IX cnt_2067__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12986), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i7.GSR = "ENABLED";
    FD1S3IX cnt_2067__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12986), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i8.GSR = "ENABLED";
    FD1S3IX cnt_2067__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12986), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module HALL_U5
//

module HALL_U5 (clk_1mhz, \speed_m1[0] , hallsense_m1, clkout_c_enable_219, 
            clkout_c_enable_244, H_A_m1_c, H_B_m1_c, H_C_m1_c, \speed_m1[1] , 
            \speed_m1[2] , \speed_m1[3] , \speed_m1[4] , \speed_m1[5] , 
            \speed_m1[6] , \speed_m1[7] , \speed_m1[8] , \speed_m1[9] , 
            \speed_m1[10] , \speed_m1[11] , \speed_m1[12] , \speed_m1[13] , 
            \speed_m1[14] , \speed_m1[15] , \speed_m1[16] , \speed_m1[17] , 
            \speed_m1[18] , \speed_m1[19] , n22378, GND_net);
    input clk_1mhz;
    output \speed_m1[0] ;
    output [2:0]hallsense_m1;
    input clkout_c_enable_219;
    input clkout_c_enable_244;
    input H_A_m1_c;
    input H_B_m1_c;
    input H_C_m1_c;
    output \speed_m1[1] ;
    output \speed_m1[2] ;
    output \speed_m1[3] ;
    output \speed_m1[4] ;
    output \speed_m1[5] ;
    output \speed_m1[6] ;
    output \speed_m1[7] ;
    output \speed_m1[8] ;
    output \speed_m1[9] ;
    output \speed_m1[10] ;
    output \speed_m1[11] ;
    output \speed_m1[12] ;
    output \speed_m1[13] ;
    output \speed_m1[14] ;
    output \speed_m1[15] ;
    output \speed_m1[16] ;
    output \speed_m1[17] ;
    output \speed_m1[18] ;
    output \speed_m1[19] ;
    input n22378;
    input GND_net;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(62[10:22])
    
    wire stable_counting, n19059;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_lat;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_104, n4299;
    wire [19:0]n7;
    
    wire hall1_old, hall1_lat, hall2_old, hall2_lat, hall3_old, n21840, 
        n21846, stable_counting_N_1746, n20145;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(60[10:15])
    
    wire n10, n25_adj_1921, n21832, n21853, n20142;
    wire [6:0]n83;
    
    wire n20397, n12, stable_counting_N_1758, n20141, n20146, n21852, 
        n20143, n20144, n95, n21872, n21827, n13_adj_1924, n22_adj_1925, 
        n18_adj_1926, n20_adj_1927, n14_adj_1928, n20371, n20413, 
        n12_adj_1929, n20403, n20251, n20367, n20307, n4, n21904, 
        n18723, n18722, n18721, n18720, n18719, n18718, n18717, 
        n18716, n18715, n18714;
    
    FD1P3AX stable_count__i0 (.D(n19059), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n7[6]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n7[5]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n7[4]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n7[3]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i2 (.D(n7[2]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m1_c), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m1_c), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[5]), .B(n21840), .C(n21846), 
         .D(stable_counting_N_1746), .Z(n20145)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0006;
    FD1P3AX hall3_lat_59 (.D(H_C_m1_c), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    LUT4 i5_3_lut_rep_412 (.A(count[13]), .B(n10), .C(n25_adj_1921), .Z(n21832)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut_rep_412.init = 16'hfefe;
    LUT4 i18281_2_lut_2_lut_4_lut (.A(count[13]), .B(n10), .C(n25_adj_1921), 
         .D(n21846), .Z(clk_1mhz_enable_104)) /* synthesis lut_function=(A (D)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i18281_2_lut_2_lut_4_lut.init = 16'hff01;
    LUT4 i1_2_lut_3_lut_4_lut_adj_178 (.A(stable_count[4]), .B(n21853), 
         .C(n21846), .D(stable_counting_N_1746), .Z(n20142)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i1_2_lut_3_lut_4_lut_adj_178.init = 16'h0006;
    LUT4 i2347_3_lut_4_lut (.A(stable_count[4]), .B(n21853), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n83[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2347_3_lut_4_lut.init = 16'h7f80;
    LUT4 i7_4_lut (.A(n20397), .B(stable_count[6]), .C(n12), .D(stable_count[2]), 
         .Z(stable_counting_N_1758)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[7:23])
    defparam i7_4_lut.init = 16'h0010;
    LUT4 i2191_2_lut_rep_426 (.A(stable_counting), .B(stable_counting_N_1758), 
         .Z(n21846)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i2191_2_lut_rep_426.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_179 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n83[6]), .D(stable_counting_N_1746), .Z(n20141)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_179.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_180 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n83[1]), .D(stable_counting_N_1746), .Z(n20146)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_180.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_181 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21852), .D(stable_counting_N_1746), .Z(n20143)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_181.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_182 (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n83[2]), .D(stable_counting_N_1746), .Z(n20144)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_182.init = 16'h0070;
    LUT4 i18284_3_lut_4_lut (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(stable_counting_N_1746), .D(stable_count[0]), .Z(n19059)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i18284_3_lut_4_lut.init = 16'h0007;
    LUT4 i17571_4_lut (.A(stable_count[3]), .B(stable_count[4]), .C(stable_count[1]), 
         .D(stable_count[5]), .Z(n20397)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17571_4_lut.init = 16'hfffe;
    FD1P3IX speedt__i1 (.D(n7[1]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    LUT4 i4_4_lut (.A(stable_count[0]), .B(n95), .C(hall2_lat), .D(hall2_old), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[7:23])
    defparam i4_4_lut.init = 16'h8008;
    LUT4 mux_28_i2_4_lut (.A(n7[1]), .B(speedt[1]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hac0a;
    LUT4 i1_4_lut (.A(hall3_lat), .B(hall1_lat), .C(hall3_old), .D(hall1_old), 
         .Z(n95)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[7:23])
    defparam i1_4_lut.init = 16'h8421;
    LUT4 mux_28_i3_4_lut (.A(n7[2]), .B(speedt[2]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hac0a;
    LUT4 mux_28_i4_4_lut (.A(n7[3]), .B(speedt[3]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hac0a;
    LUT4 mux_28_i5_4_lut (.A(n7[4]), .B(speedt[4]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hac0a;
    LUT4 mux_28_i6_4_lut (.A(n7[5]), .B(speedt[5]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hac0a;
    LUT4 mux_28_i7_4_lut (.A(n7[6]), .B(speedt[6]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hac0a;
    LUT4 mux_28_i8_4_lut (.A(n7[7]), .B(speedt[7]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hac0a;
    LUT4 mux_28_i9_4_lut (.A(n7[8]), .B(speedt[8]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hac0a;
    LUT4 mux_28_i10_4_lut (.A(n7[9]), .B(speedt[9]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hac0a;
    LUT4 mux_28_i11_4_lut (.A(n7[10]), .B(speedt[10]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hac0a;
    LUT4 mux_28_i12_4_lut (.A(n7[11]), .B(speedt[11]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hac0a;
    LUT4 mux_28_i13_4_lut (.A(n7[12]), .B(speedt[12]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hac0a;
    LUT4 mux_28_i14_4_lut (.A(n7[13]), .B(speedt[13]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hac0a;
    LUT4 mux_28_i15_4_lut (.A(n7[14]), .B(speedt[14]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hac0a;
    LUT4 mux_28_i16_4_lut (.A(n7[15]), .B(speedt[15]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hac0a;
    LUT4 mux_28_i17_4_lut (.A(n7[16]), .B(speedt[16]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hac0a;
    LUT4 mux_28_i18_4_lut (.A(n7[17]), .B(speedt[17]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hac0a;
    LUT4 mux_28_i19_4_lut (.A(n7[18]), .B(speedt[18]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hac0a;
    LUT4 mux_28_i20_4_lut (.A(n7[19]), .B(speedt[19]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hac0a;
    LUT4 i2340_2_lut_rep_407_3_lut_4_lut (.A(stable_count[3]), .B(n21872), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21827)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2340_2_lut_rep_407_3_lut_4_lut.init = 16'h78f0;
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 mux_28_i1_4_lut (.A(n7[0]), .B(speedt[0]), .C(stable_counting_N_1758), 
         .D(n21832), .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hac0a;
    LUT4 i4_4_lut_adj_183 (.A(count[11]), .B(count[6]), .C(n13_adj_1924), 
         .D(count[7]), .Z(n10)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i4_4_lut_adj_183.init = 16'hffef;
    LUT4 i11_4_lut (.A(count[9]), .B(n22_adj_1925), .C(n18_adj_1926), 
         .D(count[4]), .Z(n13_adj_1924)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i11_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(count[5]), .B(n20_adj_1927), .C(n14_adj_1928), 
         .D(count[16]), .Z(n22_adj_1925)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i10_4_lut.init = 16'h8000;
    LUT4 i6_3_lut (.A(count[1]), .B(count[15]), .C(count[0]), .Z(n18_adj_1926)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i6_3_lut.init = 16'h0202;
    LUT4 i8_4_lut (.A(count[2]), .B(count[3]), .C(count[19]), .D(count[17]), 
         .Z(n20_adj_1927)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i2_2_lut (.A(count[18]), .B(count[14]), .Z(n14_adj_1928)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i2_3_lut (.A(count[8]), .B(count[10]), .C(count[12]), .Z(n25_adj_1921)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    FD1S3IX count__i1 (.D(n7[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n7[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n7[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n7[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n7[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n7[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n7[7]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n7[8]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n7[9]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n7[10]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n7[11]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n7[12]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n7[13]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n7[14]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n7[15]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n7[16]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n7[17]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n7[18]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n7[19]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n7[19]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n7[18]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n7[17]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i0 (.D(n7[0]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(n7[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22378), .SP(stable_counting_N_1746), 
            .CD(n20371), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3AX stable_count__i1 (.D(n20146), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3AX stable_count__i2 (.D(n20144), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n7[16]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n7[15]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n7[14]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n7[13]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n7[12]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n7[11]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n7[10]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n7[9]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3AX stable_count__i3 (.D(n20143), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    LUT4 i6_4_lut (.A(n20413), .B(n12_adj_1929), .C(stable_counting), 
         .D(n83[1]), .Z(n4299)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i6_4_lut.init = 16'h4000;
    LUT4 i17587_4_lut (.A(count[11]), .B(n20403), .C(n20251), .D(count[7]), 
         .Z(n20413)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17587_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut (.A(stable_count[0]), .B(n13_adj_1924), .C(stable_counting_N_1746), 
         .D(clk_1mhz_enable_104), .Z(n12_adj_1929)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i5_4_lut.init = 16'h0800;
    LUT4 i17577_4_lut (.A(stable_counting_N_1746), .B(n83[2]), .C(n20367), 
         .D(n20307), .Z(n20403)) /* synthesis lut_function=(A (D)+!A (B+(C+(D)))) */ ;
    defparam i17577_4_lut.init = 16'hff54;
    LUT4 i17427_2_lut (.A(count[13]), .B(count[6]), .Z(n20251)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17427_2_lut.init = 16'heeee;
    LUT4 i17483_4_lut (.A(n25_adj_1921), .B(stable_counting_N_1746), .C(n21827), 
         .D(n83[6]), .Z(n20307)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;
    defparam i17483_4_lut.init = 16'hbbba;
    LUT4 i2312_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n83[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2312_2_lut.init = 16'h6666;
    LUT4 i2_3_lut_adj_184 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(92[7:87])
    defparam i2_3_lut_adj_184.init = 16'hdede;
    LUT4 i1_4_lut_adj_185 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(92[7:87])
    defparam i1_4_lut_adj_185.init = 16'h7bde;
    LUT4 i17545_3_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(stable_counting_N_1758), .Z(n20371)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i17545_3_lut.init = 16'hc8c8;
    LUT4 i2335_2_lut_rep_420_3_lut_4_lut (.A(stable_count[2]), .B(n21904), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21840)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2335_2_lut_rep_420_3_lut_4_lut.init = 16'h8000;
    LUT4 i17425_2_lut_3_lut_4_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21904), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n20367)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i17425_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h7ff8;
    FD1P3AX stable_count__i4 (.D(n20142), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3AX stable_count__i5 (.D(n20145), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3AX stable_count__i6 (.D(n20141), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n7[8]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n7[7]), .SP(clk_1mhz_enable_104), .CD(n4299), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18723), 
          .S0(n7[19]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18722), .COUT(n18723), .S0(n7[17]), .S1(n7[18]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18721), .COUT(n18722), .S0(n7[15]), .S1(n7[16]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18720), .COUT(n18721), .S0(n7[13]), .S1(n7[14]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18719), .COUT(n18720), .S0(n7[11]), .S1(n7[12]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18718), .COUT(n18719), .S0(n7[9]), .S1(n7[10]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18717), 
          .COUT(n18718), .S0(n7[7]), .S1(n7[8]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18716), 
          .COUT(n18717), .S0(n7[5]), .S1(n7[6]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18715), 
          .COUT(n18716), .S0(n7[3]), .S1(n7[4]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18714), 
          .COUT(n18715), .S0(n7[1]), .S1(n7[2]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18714), 
          .S1(n7[0]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i2314_2_lut_rep_484 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21904)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2314_2_lut_rep_484.init = 16'h8888;
    LUT4 i2321_2_lut_rep_452_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21872)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2321_2_lut_rep_452_3_lut.init = 16'h8080;
    LUT4 i2319_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n83[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2319_2_lut_3_lut.init = 16'h7878;
    LUT4 i2326_2_lut_rep_432_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21852)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2326_2_lut_rep_432_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2328_2_lut_rep_433_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21853)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2328_2_lut_rep_433_3_lut_4_lut.init = 16'h8000;
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U1
//

module PWMGENERATOR_U1 (GND_net, PWM_m2, pwm_clk, free_m2, clkout_c_enable_219, 
            PWMdut_m2, hallsense_m2, n21911, enable_m2, n2964, n21913, 
            n2928);
    input GND_net;
    output PWM_m2;
    input pwm_clk;
    output free_m2;
    input clkout_c_enable_219;
    input [9:0]PWMdut_m2;
    input [2:0]hallsense_m2;
    output n21911;
    input enable_m2;
    output n2964;
    output n21913;
    output n2928;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(88[9:16])
    
    wire n18815;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(41[10:13])
    wire [9:0]n45;
    
    wire PWM_N_1805, n18814, free_N_1817, n18813, n10, n7, n10_adj_1919, 
        n10966, n9, n18812, n18811, n3662, n17, n16, n12987, 
        n18795, n18794, n18793, n18792, n18791, n14, n10_adj_1920;
    
    CCU2D cnt_2066_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18815), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2066_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_11.INJECT1_1 = "NO";
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m2)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=318, LSE_RLINE=318 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    CCU2D cnt_2066_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18814), 
          .COUT(n18815), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_9.INJECT1_1 = "NO";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_219), .CK(pwm_clk), 
            .Q(free_m2));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    CCU2D cnt_2066_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18813), 
          .COUT(n18814), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_7.INJECT1_1 = "NO";
    LUT4 i2_3_lut (.A(PWMdut_m2[5]), .B(PWMdut_m2[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_1919), .B(PWMdut_m2[9]), .C(PWMdut_m2[8]), 
         .D(PWMdut_m2[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2263_3_lut (.A(n10966), .B(PWMdut_m2[4]), .C(PWMdut_m2[3]), 
         .Z(n10_adj_1919)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2263_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D cnt_2066_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18812), 
          .COUT(n18813), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2066_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18811), 
          .COUT(n18812), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2066_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18811), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2066_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2066_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_1.INJECT1_1 = "NO";
    LUT4 i1794_1_lut (.A(n3662), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1794_1_lut.init = 16'h5555;
    LUT4 i18303_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n12987)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(73[6:16])
    defparam i18303_4_lut.init = 16'h0400;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    FD1S3IX cnt_2066__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12987), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i0.GSR = "ENABLED";
    LUT4 i6_4_lut (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut.init = 16'hffef;
    CCU2D sub_1792_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m2[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18795), .S1(n3662));
    defparam sub_1792_add_2_11.INIT0 = 16'h5999;
    defparam sub_1792_add_2_11.INIT1 = 16'h0000;
    defparam sub_1792_add_2_11.INJECT1_0 = "NO";
    defparam sub_1792_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_9 (.A0(PWMdut_m2[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m2[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18794), 
          .COUT(n18795));
    defparam sub_1792_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1792_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1792_add_2_9.INJECT1_0 = "NO";
    defparam sub_1792_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_7 (.A0(PWMdut_m2[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m2[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18793), 
          .COUT(n18794));
    defparam sub_1792_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1792_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1792_add_2_7.INJECT1_0 = "NO";
    defparam sub_1792_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_5 (.A0(PWMdut_m2[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m2[4]), .C1(n9), .D1(n10), .CIN(n18792), 
          .COUT(n18793));
    defparam sub_1792_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1792_add_2_5.INIT1 = 16'h5999;
    defparam sub_1792_add_2_5.INJECT1_0 = "NO";
    defparam sub_1792_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m2[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m2[2]), .C1(n9), .D1(n10), .CIN(n18791), 
          .COUT(n18792));
    defparam sub_1792_add_2_3.INIT0 = 16'h5999;
    defparam sub_1792_add_2_3.INIT1 = 16'h5999;
    defparam sub_1792_add_2_3.INJECT1_0 = "NO";
    defparam sub_1792_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m2[0]), .C1(n9), .D1(n10), 
          .COUT(n18791));
    defparam sub_1792_add_2_1.INIT0 = 16'h0000;
    defparam sub_1792_add_2_1.INIT1 = 16'h5999;
    defparam sub_1792_add_2_1.INJECT1_0 = "NO";
    defparam sub_1792_add_2_1.INJECT1_1 = "NO";
    LUT4 i18257_4_lut (.A(PWMdut_m2[5]), .B(n14), .C(n10_adj_1920), .D(PWMdut_m2[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i18257_4_lut.init = 16'h0001;
    LUT4 i6_4_lut_adj_176 (.A(PWMdut_m2[9]), .B(PWMdut_m2[3]), .C(PWMdut_m2[4]), 
         .D(n10966), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut_adj_176.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[7]), .Z(n10_adj_1920)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_177 (.A(PWMdut_m2[2]), .B(PWMdut_m2[1]), .C(PWMdut_m2[0]), 
         .Z(n10966)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_177.init = 16'hfefe;
    LUT4 i1538_3_lut_rep_491 (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .Z(n21911)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1538_3_lut_rep_491.init = 16'h1414;
    LUT4 i18341_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .D(enable_m2), .Z(n2964)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18341_2_lut_4_lut.init = 16'hebff;
    LUT4 i1508_3_lut_rep_493 (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .Z(n21913)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1508_3_lut_rep_493.init = 16'h1414;
    LUT4 i18338_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .D(enable_m2), .Z(n2928)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18338_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2066__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12987), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i1.GSR = "ENABLED";
    FD1S3IX cnt_2066__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12987), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i2.GSR = "ENABLED";
    FD1S3IX cnt_2066__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12987), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i3.GSR = "ENABLED";
    FD1S3IX cnt_2066__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12987), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i4.GSR = "ENABLED";
    FD1S3IX cnt_2066__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12987), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i5.GSR = "ENABLED";
    FD1S3IX cnt_2066__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12987), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i6.GSR = "ENABLED";
    FD1S3IX cnt_2066__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12987), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i7.GSR = "ENABLED";
    FD1S3IX cnt_2066__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12987), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i8.GSR = "ENABLED";
    FD1S3IX cnt_2066__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12987), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U2
//

module PWMGENERATOR_U2 (GND_net, PWM_m1, pwm_clk, free_m1, clkout_c_enable_244, 
            PWMdut_m1, hallsense_m1, n21920, enable_m1, n2798, n2834, 
            n21918);
    input GND_net;
    output PWM_m1;
    input pwm_clk;
    output free_m1;
    input clkout_c_enable_244;
    input [9:0]PWMdut_m1;
    input [2:0]hallsense_m1;
    output n21920;
    input enable_m1;
    output n2798;
    output n2834;
    output n21918;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(88[9:16])
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(41[10:13])
    wire [9:0]n45;
    
    wire n18816, PWM_N_1805, free_N_1817, n10, n7, n10_adj_1917, 
        n10964, n9, n3649, n20407, n6, n12988, n20381, n18800, 
        n18799, n18798, n18797, n18796, n14, n10_adj_1918, n18820, 
        n18819, n18818, n18817;
    
    CCU2D cnt_2065_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18816), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2065_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2065_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_1.INJECT1_1 = "NO";
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=308, LSE_RLINE=308 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_244), .CK(pwm_clk), 
            .Q(free_m1));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(PWMdut_m1[5]), .B(PWMdut_m1[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_1917), .B(PWMdut_m1[9]), .C(PWMdut_m1[8]), 
         .D(PWMdut_m1[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2266_3_lut (.A(n10964), .B(PWMdut_m1[4]), .C(PWMdut_m1[3]), 
         .Z(n10_adj_1917)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2266_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1792_1_lut (.A(n3649), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1792_1_lut.init = 16'h5555;
    LUT4 i18306_4_lut (.A(cnt[0]), .B(n20407), .C(cnt[2]), .D(n6), .Z(n12988)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(73[6:16])
    defparam i18306_4_lut.init = 16'h0004;
    LUT4 i17581_3_lut (.A(cnt[7]), .B(n20381), .C(cnt[3]), .Z(n20407)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17581_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i17555_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n20381)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17555_4_lut.init = 16'h8000;
    FD1S3IX cnt_2065__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12988), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i0.GSR = "ENABLED";
    CCU2D sub_1790_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m1[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18800), .S1(n3649));
    defparam sub_1790_add_2_11.INIT0 = 16'h5999;
    defparam sub_1790_add_2_11.INIT1 = 16'h0000;
    defparam sub_1790_add_2_11.INJECT1_0 = "NO";
    defparam sub_1790_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_9 (.A0(PWMdut_m1[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m1[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18799), 
          .COUT(n18800));
    defparam sub_1790_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1790_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1790_add_2_9.INJECT1_0 = "NO";
    defparam sub_1790_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_7 (.A0(PWMdut_m1[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m1[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18798), 
          .COUT(n18799));
    defparam sub_1790_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1790_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1790_add_2_7.INJECT1_0 = "NO";
    defparam sub_1790_add_2_7.INJECT1_1 = "NO";
    LUT4 i1416_3_lut_rep_500 (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .Z(n21920)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1416_3_lut_rep_500.init = 16'h1414;
    CCU2D sub_1790_add_2_5 (.A0(PWMdut_m1[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m1[4]), .C1(n9), .D1(n10), .CIN(n18797), 
          .COUT(n18798));
    defparam sub_1790_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1790_add_2_5.INIT1 = 16'h5999;
    defparam sub_1790_add_2_5.INJECT1_0 = "NO";
    defparam sub_1790_add_2_5.INJECT1_1 = "NO";
    LUT4 i18328_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .D(enable_m1), .Z(n2798)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18328_2_lut_4_lut.init = 16'hebff;
    CCU2D sub_1790_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m1[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m1[2]), .C1(n9), .D1(n10), .CIN(n18796), 
          .COUT(n18797));
    defparam sub_1790_add_2_3.INIT0 = 16'h5999;
    defparam sub_1790_add_2_3.INIT1 = 16'h5999;
    defparam sub_1790_add_2_3.INJECT1_0 = "NO";
    defparam sub_1790_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m1[0]), .C1(n9), .D1(n10), 
          .COUT(n18796));
    defparam sub_1790_add_2_1.INIT0 = 16'h0000;
    defparam sub_1790_add_2_1.INIT1 = 16'h5999;
    defparam sub_1790_add_2_1.INJECT1_0 = "NO";
    defparam sub_1790_add_2_1.INJECT1_1 = "NO";
    LUT4 i18260_4_lut (.A(PWMdut_m1[5]), .B(n14), .C(n10_adj_1918), .D(PWMdut_m1[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i18260_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m1[9]), .B(PWMdut_m1[3]), .C(PWMdut_m1[4]), 
         .D(n10964), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[7]), .Z(n10_adj_1918)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_175 (.A(PWMdut_m1[2]), .B(PWMdut_m1[1]), .C(PWMdut_m1[0]), 
         .Z(n10964)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_175.init = 16'hfefe;
    LUT4 i18331_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .D(enable_m1), .Z(n2834)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i18331_2_lut_4_lut.init = 16'hebff;
    LUT4 i1446_3_lut_rep_498 (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .Z(n21918)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(52[2] 76[9])
    defparam i1446_3_lut_rep_498.init = 16'h1414;
    FD1S3IX cnt_2065__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12988), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i1.GSR = "ENABLED";
    FD1S3IX cnt_2065__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12988), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i2.GSR = "ENABLED";
    FD1S3IX cnt_2065__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12988), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i3.GSR = "ENABLED";
    FD1S3IX cnt_2065__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12988), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i4.GSR = "ENABLED";
    FD1S3IX cnt_2065__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12988), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i5.GSR = "ENABLED";
    FD1S3IX cnt_2065__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12988), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i6.GSR = "ENABLED";
    FD1S3IX cnt_2065__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12988), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i7.GSR = "ENABLED";
    FD1S3IX cnt_2065__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12988), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i8.GSR = "ENABLED";
    FD1S3IX cnt_2065__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12988), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i9.GSR = "ENABLED";
    CCU2D cnt_2065_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18820), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2065_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18819), 
          .COUT(n18820), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18818), 
          .COUT(n18819), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18817), 
          .COUT(n18818), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18816), 
          .COUT(n18817), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_3.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module HALL_U4
//

module HALL_U4 (clk_1mhz, \speed_m2[0] , hallsense_m2, clkout_c_enable_244, 
            clkout_c_enable_219, H_C_m2_c, H_B_m2_c, H_A_m2_c, \speed_m2[1] , 
            \speed_m2[2] , \speed_m2[3] , \speed_m2[4] , \speed_m2[5] , 
            \speed_m2[6] , \speed_m2[7] , \speed_m2[8] , \speed_m2[9] , 
            \speed_m2[10] , \speed_m2[11] , \speed_m2[12] , \speed_m2[13] , 
            \speed_m2[14] , \speed_m2[15] , \speed_m2[16] , \speed_m2[17] , 
            \speed_m2[18] , \speed_m2[19] , n22378, GND_net);
    input clk_1mhz;
    output \speed_m2[0] ;
    output [2:0]hallsense_m2;
    input clkout_c_enable_244;
    input clkout_c_enable_219;
    input H_C_m2_c;
    input H_B_m2_c;
    input H_A_m2_c;
    output \speed_m2[1] ;
    output \speed_m2[2] ;
    output \speed_m2[3] ;
    output \speed_m2[4] ;
    output \speed_m2[5] ;
    output \speed_m2[6] ;
    output \speed_m2[7] ;
    output \speed_m2[8] ;
    output \speed_m2[9] ;
    output \speed_m2[10] ;
    output \speed_m2[11] ;
    output \speed_m2[12] ;
    output \speed_m2[13] ;
    output \speed_m2[14] ;
    output \speed_m2[15] ;
    output \speed_m2[16] ;
    output \speed_m2[17] ;
    output \speed_m2[18] ;
    output \speed_m2[19] ;
    input n22378;
    input GND_net;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(62[10:22])
    
    wire stable_counting, n19064;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_lat, hall3_old, hall1_old, hall1_lat, hall2_lat;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_83, n4334;
    wire [19:0]n1;
    
    wire hall2_old;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(60[10:15])
    
    wire n16, n12, n21829, n21844;
    wire [6:0]n83;
    
    wire n20223, n21861, n20148, n13, n19132, n21881, stable_counting_N_1746, 
        n7, n20153, n20149, n20150, n20151, n20152, n21880, n21833, 
        n20319, n20337, n19_adj_1909, n20345, n20327, n20287, n21876, 
        n10_adj_1910, n5216, n4, n20214, n15_adj_1911, n21921, n21845, 
        n18733, n18732, n18731, n18730, n18729, n18728, n18727, 
        n18726, n18725, n18724, n18_adj_1912, n14_adj_1913, n12_adj_1914, 
        n20_adj_1915, n17_adj_1916, n20339;
    
    FD1P3AX stable_count__i0 (.D(n19064), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m2_c), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m2_c), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3IX speedt__i0 (.D(n1[0]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 i8_4_lut_rep_409 (.A(count[7]), .B(n16), .C(n12), .D(count[15]), 
         .Z(n21829)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_4_lut_rep_409.init = 16'hfffe;
    LUT4 i17399_3_lut_4_lut (.A(stable_count[5]), .B(n21844), .C(n83[6]), 
         .D(n83[3]), .Z(n20223)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i17399_3_lut_4_lut.init = 16'hfff6;
    LUT4 i2397_3_lut_4_lut (.A(stable_count[4]), .B(n21861), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n83[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2397_3_lut_4_lut.init = 16'h7f80;
    FD1P3AX hall1_lat_57 (.D(H_A_m2_c), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX stable_count__i6 (.D(n20148), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    LUT4 mux_28_i2_4_lut (.A(n1[1]), .B(speedt[1]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i3_4_lut (.A(n1[2]), .B(speedt[2]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i4_4_lut (.A(n1[3]), .B(speedt[3]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i5_4_lut (.A(n1[4]), .B(speedt[4]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i6_4_lut (.A(n1[5]), .B(speedt[5]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i7_4_lut (.A(n1[6]), .B(speedt[6]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i8_4_lut (.A(n1[7]), .B(speedt[7]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i9_4_lut (.A(n1[8]), .B(speedt[8]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i10_4_lut (.A(n1[9]), .B(speedt[9]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i11_4_lut (.A(n1[10]), .B(speedt[10]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i12_4_lut (.A(n1[11]), .B(speedt[11]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i13_4_lut (.A(n1[12]), .B(speedt[12]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i14_4_lut (.A(n1[13]), .B(speedt[13]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i15_4_lut (.A(n1[14]), .B(speedt[14]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i16_4_lut (.A(n1[15]), .B(speedt[15]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i17_4_lut (.A(n1[16]), .B(speedt[16]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i18_4_lut (.A(n1[17]), .B(speedt[17]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i19_4_lut (.A(n1[18]), .B(speedt[18]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i20_4_lut (.A(n1[19]), .B(speedt[19]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hcaa0;
    LUT4 i3_4_lut (.A(n19132), .B(n21881), .C(stable_counting_N_1746), 
         .D(n83[1]), .Z(n13)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[7:23])
    defparam i3_4_lut.init = 16'hfeff;
    LUT4 i4_4_lut (.A(n7), .B(n83[6]), .C(stable_count[0]), .D(n83[3]), 
         .Z(n19132)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[7:23])
    defparam i4_4_lut.init = 16'hffef;
    LUT4 i2362_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n83[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2362_2_lut.init = 16'h6666;
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n1[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n1[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n1[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n1[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n1[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n1[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n1[7]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n1[8]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n1[9]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n1[10]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n1[11]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n1[12]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n1[13]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n1[14]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n1[15]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n1[16]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n1[17]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n1[18]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n1[19]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3AX stable_count__i5 (.D(n20153), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3AX stable_count__i4 (.D(n20149), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3AX stable_count__i3 (.D(n20150), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3AX stable_count__i2 (.D(n20151), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3AX stable_count__i1 (.D(n20152), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    LUT4 i2390_2_lut_rep_413_3_lut_4_lut (.A(stable_count[3]), .B(n21880), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21833)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2390_2_lut_rep_413_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2_2_lut_3_lut_4_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21880), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n7)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h7ff8;
    LUT4 i17494_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21880), .C(n21881), 
         .D(stable_count[4]), .Z(n20319)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (C+(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i17494_2_lut_3_lut_4_lut.init = 16'hf7f8;
    LUT4 i18287_2_lut_3_lut_3_lut_4_lut (.A(stable_count[0]), .B(stable_counting_N_1746), 
         .C(stable_counting), .D(n13), .Z(n19064)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i18287_2_lut_3_lut_3_lut_4_lut.init = 16'h1101;
    LUT4 i8_3_lut_4_lut (.A(stable_count[0]), .B(stable_counting_N_1746), 
         .C(count[12]), .D(n20337), .Z(n19_adj_1909)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i8_3_lut_4_lut.init = 16'h000e;
    LUT4 mux_28_i1_4_lut (.A(n1[0]), .B(speedt[0]), .C(n13), .D(n21829), 
         .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hcaa0;
    LUT4 i7_4_lut (.A(n20337), .B(n20345), .C(n20327), .D(n20287), .Z(n16)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i7_4_lut.init = 16'hfbff;
    LUT4 i3_2_lut (.A(count[6]), .B(count[12]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i17520_4_lut (.A(count[13]), .B(count[1]), .C(n21876), .D(count[2]), 
         .Z(n20345)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i17520_4_lut.init = 16'h4000;
    LUT4 i17463_3_lut (.A(count[4]), .B(count[17]), .C(count[3]), .Z(n20287)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17463_3_lut.init = 16'h8080;
    LUT4 i4_4_lut_adj_166 (.A(count[9]), .B(count[5]), .C(count[19]), 
         .D(count[16]), .Z(n10_adj_1910)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut_adj_166.init = 16'h8000;
    LUT4 i17512_2_lut (.A(count[0]), .B(count[10]), .Z(n20337)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17512_2_lut.init = 16'heeee;
    LUT4 i17502_2_lut (.A(count[8]), .B(count[11]), .Z(n20327)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17502_2_lut.init = 16'heeee;
    FD1P3IX speedt__i1 (.D(n1[1]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(n1[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_83), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22378), .SP(stable_counting_N_1746), 
            .CD(n5216), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3IX speedt__i2 (.D(n1[2]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n1[3]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n1[4]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n1[5]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n1[6]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n1[7]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n1[8]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n1[9]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n1[10]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n1[11]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n1[12]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n1[13]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n1[14]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n1[15]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n1[16]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n1[17]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n1[18]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n1[19]), .SP(clk_1mhz_enable_83), .CD(n4334), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(hall2_old), .B(hall1_old), .C(hall2_lat), .D(hall1_lat), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(92[7:87])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i18268_4_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(n83[1]), .D(n20214), .Z(n5216)) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(97[3] 113[10])
    defparam i18268_4_lut.init = 16'h88c8;
    LUT4 i5_3_lut_rep_456 (.A(count[18]), .B(n10_adj_1910), .C(count[14]), 
         .Z(n21876)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut_rep_456.init = 16'h8080;
    LUT4 i5_2_lut_4_lut (.A(count[18]), .B(n10_adj_1910), .C(count[14]), 
         .D(n83[1]), .Z(n15_adj_1911)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_2_lut_4_lut.init = 16'h8000;
    LUT4 i2385_2_lut_rep_424_3_lut_4_lut (.A(stable_count[2]), .B(n21921), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21844)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2385_2_lut_rep_424_3_lut_4_lut.init = 16'h8000;
    LUT4 i2383_2_lut_rep_425_3_lut_4_lut (.A(stable_count[2]), .B(n21921), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21845)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2383_2_lut_rep_425_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2_3_lut_rep_462 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_462.init = 16'hdede;
    LUT4 i2364_2_lut_rep_501 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21921)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2364_2_lut_rep_501.init = 16'h8888;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18733), 
          .S0(n1[19]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18732), .COUT(n18733), .S0(n1[17]), .S1(n1[18]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18731), .COUT(n18732), .S0(n1[15]), .S1(n1[16]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18730), .COUT(n18731), .S0(n1[13]), .S1(n1[14]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18729), .COUT(n18730), .S0(n1[11]), .S1(n1[12]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18728), .COUT(n18729), .S0(n1[9]), .S1(n1[10]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18727), 
          .COUT(n18728), .S0(n1[7]), .S1(n1[8]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18726), 
          .COUT(n18727), .S0(n1[5]), .S1(n1[6]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18725), 
          .COUT(n18726), .S0(n1[3]), .S1(n1[4]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18724), 
          .COUT(n18725), .S0(n1[1]), .S1(n1[2]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18724), 
          .S1(n1[0]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i2371_2_lut_rep_460_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21880)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2371_2_lut_rep_460_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_counting), .B(n13), .C(n83[1]), 
         .D(stable_counting_N_1746), .Z(n20152)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h00d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_167 (.A(stable_counting), .B(n13), .C(n21845), 
         .D(stable_counting_N_1746), .Z(n20149)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_167.init = 16'h00d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_168 (.A(stable_counting), .B(n13), .C(n21833), 
         .D(stable_counting_N_1746), .Z(n20153)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_168.init = 16'h00d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_169 (.A(stable_counting), .B(n13), .C(n83[6]), 
         .D(stable_counting_N_1746), .Z(n20148)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_169.init = 16'h00d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_170 (.A(stable_counting), .B(n13), .C(n83[3]), 
         .D(stable_counting_N_1746), .Z(n20150)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_170.init = 16'h00d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_171 (.A(stable_counting), .B(n13), .C(n21881), 
         .D(stable_counting_N_1746), .Z(n20151)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_171.init = 16'h00d0;
    LUT4 i9_4_lut (.A(count[4]), .B(n18_adj_1912), .C(n14_adj_1913), .D(count[3]), 
         .Z(n4334)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i8_4_lut (.A(n15_adj_1911), .B(stable_counting), .C(n12_adj_1914), 
         .D(stable_counting_N_1746), .Z(n18_adj_1912)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i8_4_lut.init = 16'h0080;
    LUT4 i4_4_lut_adj_172 (.A(count[17]), .B(clk_1mhz_enable_83), .C(n19_adj_1909), 
         .D(n20_adj_1915), .Z(n14_adj_1913)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut_adj_172.init = 16'h8000;
    LUT4 i2_2_lut (.A(count[2]), .B(count[1]), .Z(n12_adj_1914)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i9_4_lut_adj_173 (.A(n17_adj_1916), .B(count[6]), .C(n20339), 
         .D(count[15]), .Z(n20_adj_1915)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i9_4_lut_adj_173.init = 16'h0002;
    LUT4 i6_4_lut (.A(n20223), .B(n20327), .C(stable_counting_N_1746), 
         .D(n20319), .Z(n17_adj_1916)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i6_4_lut.init = 16'h3031;
    LUT4 i17514_2_lut (.A(count[13]), .B(count[7]), .Z(n20339)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17514_2_lut.init = 16'heeee;
    LUT4 i18276_2_lut_3_lut_3_lut (.A(n21829), .B(n13), .C(stable_counting), 
         .Z(clk_1mhz_enable_83)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i18276_2_lut_3_lut_3_lut.init = 16'h7575;
    LUT4 i2378_2_lut_rep_441_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21861)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2378_2_lut_rep_441_3_lut_4_lut.init = 16'h8000;
    LUT4 i2376_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n83[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2376_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2369_2_lut_rep_461_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21881)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2369_2_lut_rep_461_3_lut.init = 16'h7878;
    LUT4 i1_2_lut_3_lut_4_lut_adj_174 (.A(stable_count[1]), .B(stable_count[0]), 
         .C(n19132), .D(stable_count[2]), .Z(n20214)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (C+(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i1_2_lut_3_lut_4_lut_adj_174.init = 16'hf7f8;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module SPI
//

module SPI (MISO_N_624, clkout_c, enable_m4, clkout_c_enable_219, speed_set_m3, 
            HALL_A_OUT_c_c, clkout_c_enable_244, HALL_B_OUT_c_c, enable_m1, 
            free_m1, hallsense_m1, n20053, enable_m2, n21864, enable_m3, 
            HALL_C_OUT_c_c, n21865, dir_m1, n2786, n2822, hallsense_m2, 
            dir_m2, n2916, n2952, speed_set_m4, hallsense_m3, n21907, 
            dir_m3, n3046, n3082, speed_set_m2, n22383, rst, \send_buffer[94] , 
            \send_buffer_95__N_346[94] , hallsense_m4, dir_m4, n3176, 
            n3212, GND_net, speed_set_m1, \speed_m1[19] , \speed_m2[1] , 
            \speed_m2[2] , \speed_m3[19] , \speed_m2[3] , \speed_m2[0] , 
            \speed_m2[4] , \speed_m2[5] , \speed_m2[6] , \speed_m2[7] , 
            \speed_m2[8] , \speed_m2[9] , \speed_m2[10] , \speed_m2[11] , 
            \speed_m2[12] , \speed_m2[13] , \speed_m2[14] , \speed_m2[15] , 
            \speed_m2[16] , \speed_m2[17] , \speed_m4[6] , \speed_m4[5] , 
            \speed_m2[18] , \speed_m2[19] , \speed_m1[0] , \speed_m1[1] , 
            \speed_m1[2] , \speed_m1[3] , \speed_m1[4] , \speed_m1[5] , 
            \speed_m1[6] , \speed_m1[7] , \speed_m1[8] , \speed_m1[9] , 
            \speed_m1[10] , \speed_m1[11] , \speed_m1[12] , \speed_m1[13] , 
            \speed_m1[14] , \speed_m1[15] , \speed_m1[16] , \speed_m4[8] , 
            \speed_m4[7] , \speed_m1[17] , \speed_m1[18] , \speed_m4[10] , 
            \speed_m4[9] , \speed_m4[11] , \speed_m4[12] , \speed_m4[13] , 
            \speed_m4[14] , \speed_m4[15] , \speed_m4[16] , \speed_m4[17] , 
            \speed_m4[18] , \speed_m4[19] , \speed_m3[0] , \speed_m3[1] , 
            \speed_m3[2] , \speed_m3[3] , \speed_m3[4] , \speed_m3[5] , 
            \speed_m3[6] , \speed_m3[7] , \speed_m3[8] , \speed_m3[9] , 
            n4884, \speed_m3[10] , \speed_m3[11] , \speed_m3[12] , \speed_m3[13] , 
            \speed_m3[14] , \speed_m3[15] , \speed_m3[16] , \speed_m3[17] , 
            \speed_m3[18] , \speed_m4[0] , \speed_m4[1] , \speed_m4[2] , 
            \speed_m4[3] , \speed_m4[4] , free_m4, n20030, free_m2, 
            n20041);
    output MISO_N_624;
    input clkout_c;
    output enable_m4;
    input clkout_c_enable_219;
    output [20:0]speed_set_m3;
    input HALL_A_OUT_c_c;
    input clkout_c_enable_244;
    input HALL_B_OUT_c_c;
    output enable_m1;
    input free_m1;
    input [2:0]hallsense_m1;
    output n20053;
    output enable_m2;
    output n21864;
    output enable_m3;
    input HALL_C_OUT_c_c;
    output n21865;
    input dir_m1;
    output n2786;
    output n2822;
    input [2:0]hallsense_m2;
    input dir_m2;
    output n2916;
    output n2952;
    output [20:0]speed_set_m4;
    input [2:0]hallsense_m3;
    input n21907;
    input dir_m3;
    output n3046;
    output n3082;
    output [20:0]speed_set_m2;
    input n22383;
    input rst;
    output \send_buffer[94] ;
    input \send_buffer_95__N_346[94] ;
    input [2:0]hallsense_m4;
    input dir_m4;
    output n3176;
    output n3212;
    input GND_net;
    output [20:0]speed_set_m1;
    input \speed_m1[19] ;
    input \speed_m2[1] ;
    input \speed_m2[2] ;
    input \speed_m3[19] ;
    input \speed_m2[3] ;
    input \speed_m2[0] ;
    input \speed_m2[4] ;
    input \speed_m2[5] ;
    input \speed_m2[6] ;
    input \speed_m2[7] ;
    input \speed_m2[8] ;
    input \speed_m2[9] ;
    input \speed_m2[10] ;
    input \speed_m2[11] ;
    input \speed_m2[12] ;
    input \speed_m2[13] ;
    input \speed_m2[14] ;
    input \speed_m2[15] ;
    input \speed_m2[16] ;
    input \speed_m2[17] ;
    input \speed_m4[6] ;
    input \speed_m4[5] ;
    input \speed_m2[18] ;
    input \speed_m2[19] ;
    input \speed_m1[0] ;
    input \speed_m1[1] ;
    input \speed_m1[2] ;
    input \speed_m1[3] ;
    input \speed_m1[4] ;
    input \speed_m1[5] ;
    input \speed_m1[6] ;
    input \speed_m1[7] ;
    input \speed_m1[8] ;
    input \speed_m1[9] ;
    input \speed_m1[10] ;
    input \speed_m1[11] ;
    input \speed_m1[12] ;
    input \speed_m1[13] ;
    input \speed_m1[14] ;
    input \speed_m1[15] ;
    input \speed_m1[16] ;
    input \speed_m4[8] ;
    input \speed_m4[7] ;
    input \speed_m1[17] ;
    input \speed_m1[18] ;
    input \speed_m4[10] ;
    input \speed_m4[9] ;
    input \speed_m4[11] ;
    input \speed_m4[12] ;
    input \speed_m4[13] ;
    input \speed_m4[14] ;
    input \speed_m4[15] ;
    input \speed_m4[16] ;
    input \speed_m4[17] ;
    input \speed_m4[18] ;
    input \speed_m4[19] ;
    input \speed_m3[0] ;
    input \speed_m3[1] ;
    input \speed_m3[2] ;
    input \speed_m3[3] ;
    input \speed_m3[4] ;
    input \speed_m3[5] ;
    input \speed_m3[6] ;
    input \speed_m3[7] ;
    input \speed_m3[8] ;
    input \speed_m3[9] ;
    output n4884;
    input \speed_m3[10] ;
    input \speed_m3[11] ;
    input \speed_m3[12] ;
    input \speed_m3[13] ;
    input \speed_m3[14] ;
    input \speed_m3[15] ;
    input \speed_m3[16] ;
    input \speed_m3[17] ;
    input \speed_m3[18] ;
    input \speed_m4[0] ;
    input \speed_m4[1] ;
    input \speed_m4[2] ;
    input \speed_m4[3] ;
    input \speed_m4[4] ;
    input free_m4;
    output n20030;
    input free_m2;
    output n20041;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(44[2:8])
    
    wire MISO_N_670, enable_m1_N_633, enable_m4_N_649, CSold, CSlatched, 
        SCKold, SCKlatched, clkout_c_enable_245, n13012;
    wire [95:0]recv_buffer;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(68[10:21])
    wire [83:0]n169;
    
    wire clkout_c_enable_64, enable_m1_N_627, n21919, enable_m2_N_635, 
        n21887;
    wire [95:0]send_buffer;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(67[10:21])
    
    wire MISOb, n21812, enable_m3_N_642, MISO_N_625, n21889, MISOb_N_660, 
        clkout_c_enable_99;
    wire [95:0]MISOb_N_666;
    wire [95:0]send_buffer_95__N_346;
    
    wire n3480, n3456, n39, n40, n36, n28, n38, n32, n34, 
        n24, n3432, n3408, n39_adj_1874, n40_adj_1875, n36_adj_1876, 
        n28_adj_1877, n38_adj_1878, n32_adj_1879, n21912, n12992, 
        n34_adj_1880, n24_adj_1881, n13032, n21901, n21813, n18895, 
        n3336, n18894, n18893, n18892, n18891, n18890, n3312, 
        n39_adj_1882, n40_adj_1883, n18889, n36_adj_1884, n28_adj_1885, 
        n38_adj_1886, n32_adj_1887, n13052, n18888, n34_adj_1888, 
        n24_adj_1889, n18887, n18886, n18885, n18884, n22382, n18883, 
        n18882, n22381, n21863, n18881, n18880, n18879, n18971, 
        n18970, n18969, n18968, n18967, n18966, n18965, n18964, 
        n18963, n18962, n18961, n18960, n18959, n18958, n18957, 
        n18956, n18955, n18954, n18953, n18952, n18951, n18950, 
        n18949, n18948, n18947, n18946, n18945, n18944, n18943, 
        n18942, n18941, n18940, n18939, n18938, n18937, n3384, 
        n18936, n18935, n18934, n18933, n18932, n18931, n18930, 
        n3360, n18929, n18928, n18927, n18926, n18925, n18924, 
        n18923, n18922, n18921, n39_adj_1898, n40_adj_1899, n36_adj_1900, 
        n28_adj_1901, n38_adj_1902, n32_adj_1903, n34_adj_1904, n24_adj_1905;
    
    FD1S3AX MISO_124 (.D(MISO_N_670), .CK(clkout_c), .Q(MISO_N_624)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISO_124.GSR = "DISABLED";
    FD1P3AX enable_m4_112 (.D(enable_m4_N_649), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m4));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m4_112.GSR = "ENABLED";
    FD1P3AX CSold_113 (.D(CSlatched), .SP(clkout_c_enable_219), .CK(clkout_c), 
            .Q(CSold));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_113.GSR = "DISABLED";
    FD1P3AX SCKold_114 (.D(SCKlatched), .SP(clkout_c_enable_219), .CK(clkout_c), 
            .Q(SCKold));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKold_114.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i1 (.D(recv_buffer[34]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i1.GSR = "DISABLED";
    FD1P3AX CSlatched_115 (.D(HALL_A_OUT_c_c), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(CSlatched));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_115.GSR = "DISABLED";
    FD1P3AX SCKlatched_116 (.D(HALL_B_OUT_c_c), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(SCKlatched));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKlatched_116.GSR = "DISABLED";
    FD1P3AX \SPI__7_rep_4__i0  (.D(recv_buffer[13]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(n169[0]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7_rep_4__i0 .GSR = "DISABLED";
    FD1P3AX enable_m1_109 (.D(enable_m1_N_627), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m1));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m1_109.GSR = "ENABLED";
    FD1P3JX speed_set_m3_i0_i2 (.D(recv_buffer[35]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i2.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i3 (.D(recv_buffer[36]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i4 (.D(recv_buffer[37]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i4.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_499 (.A(enable_m1), .B(free_m1), .Z(n21919)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_499.init = 16'h2222;
    LUT4 i18335_3_lut_4_lut (.A(enable_m1), .B(free_m1), .C(hallsense_m1[2]), 
         .D(hallsense_m1[0]), .Z(n20053)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i18335_3_lut_4_lut.init = 16'hfddf;
    FD1P3AX enable_m2_110 (.D(enable_m2_N_635), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m2));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m2_110.GSR = "ENABLED";
    LUT4 MISOb_N_667_bdd_4_lut (.A(n21887), .B(send_buffer[1]), .C(MISOb), 
         .D(n21864), .Z(n21812)) /* synthesis lut_function=(A (B+(D))+!A !((D)+!C)) */ ;
    defparam MISOb_N_667_bdd_4_lut.init = 16'haad8;
    FD1P3AX enable_m3_111 (.D(enable_m3_N_642), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m3));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m3_111.GSR = "ENABLED";
    FD1P3AX i101_125 (.D(n21889), .SP(clkout_c_enable_219), .CK(clkout_c), 
            .Q(MISO_N_625));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i101_125.GSR = "DISABLED";
    FD1P3AX MISOb_118 (.D(MISOb_N_660), .SP(clkout_c_enable_244), .CK(clkout_c), 
            .Q(MISOb));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISOb_118.GSR = "DISABLED";
    FD1P3AX \SPI__7__i83  (.D(HALL_C_OUT_c_c), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[95]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i83 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i82  (.D(recv_buffer[95]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[94]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i82 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i81  (.D(recv_buffer[94]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[93]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i81 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i80  (.D(recv_buffer[93]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[92]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i80 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i79  (.D(recv_buffer[92]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[91]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i79 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i78  (.D(recv_buffer[91]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[90]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i78 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i77  (.D(recv_buffer[90]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[89]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i77 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i76  (.D(recv_buffer[89]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[88]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i76 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i75  (.D(recv_buffer[88]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[87]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i75 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i74  (.D(recv_buffer[87]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[86]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i74 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i73  (.D(recv_buffer[86]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[85]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i73 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i72  (.D(recv_buffer[85]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[84]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i72 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i71  (.D(recv_buffer[84]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[83]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i71 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i70  (.D(recv_buffer[83]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[82]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i70 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i69  (.D(recv_buffer[82]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[81]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i69 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i68  (.D(recv_buffer[81]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[80]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i68 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i67  (.D(recv_buffer[80]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[79]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i67 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i66  (.D(recv_buffer[79]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[78]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i66 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i65  (.D(recv_buffer[78]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[77]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i65 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i64  (.D(recv_buffer[77]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[76]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i64 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i63  (.D(recv_buffer[76]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[75]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i63 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i62  (.D(recv_buffer[75]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[74]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i62 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i61  (.D(recv_buffer[74]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[73]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i61 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i60  (.D(recv_buffer[73]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[72]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i60 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i59  (.D(recv_buffer[72]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[71]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i59 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i58  (.D(recv_buffer[71]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[70]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i58 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i57  (.D(recv_buffer[70]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[69]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i57 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i56  (.D(recv_buffer[69]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[68]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i56 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i55  (.D(recv_buffer[68]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[67]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i55 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i54  (.D(recv_buffer[67]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[66]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i54 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i53  (.D(recv_buffer[66]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[65]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i53 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i52  (.D(recv_buffer[65]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[64]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i52 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i51  (.D(recv_buffer[64]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[63]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i51 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i50  (.D(recv_buffer[63]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[62]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i50 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i49  (.D(recv_buffer[62]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[61]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i49 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i48  (.D(recv_buffer[61]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[60]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i48 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i47  (.D(recv_buffer[60]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[59]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i47 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i46  (.D(recv_buffer[59]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[58]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i46 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i45  (.D(recv_buffer[58]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[57]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i45 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i44  (.D(recv_buffer[57]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[56]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i44 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i43  (.D(recv_buffer[56]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[55]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i43 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i42  (.D(recv_buffer[55]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[54]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i42 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i41  (.D(recv_buffer[54]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[53]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i41 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i40  (.D(recv_buffer[53]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[52]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i40 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i39  (.D(recv_buffer[52]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[51]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i39 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i38  (.D(recv_buffer[51]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[50]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i38 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i37  (.D(recv_buffer[50]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[49]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i37 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i36  (.D(recv_buffer[49]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[48]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i36 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i35  (.D(recv_buffer[48]), .SP(clkout_c_enable_64), 
            .CK(clkout_c), .Q(recv_buffer[47]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i35 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i34  (.D(recv_buffer[47]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[46]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i34 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i33  (.D(recv_buffer[46]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[45]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i33 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i32  (.D(recv_buffer[45]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[44]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i32 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i31  (.D(recv_buffer[44]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[43]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i31 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i30  (.D(recv_buffer[43]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[42]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i30 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i29  (.D(recv_buffer[42]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[41]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i29 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i28  (.D(recv_buffer[41]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[40]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i28 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i27  (.D(recv_buffer[40]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[39]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i27 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i26  (.D(recv_buffer[39]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[38]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i26 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i25  (.D(recv_buffer[38]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[37]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i25 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i24  (.D(recv_buffer[37]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[36]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i24 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i23  (.D(recv_buffer[36]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[35]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i23 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i22  (.D(recv_buffer[35]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[34]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i22 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i21  (.D(recv_buffer[34]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[33]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i21 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i20  (.D(recv_buffer[33]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[32]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i20 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i19  (.D(recv_buffer[32]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[31]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i19 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i18  (.D(recv_buffer[31]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[30]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i18 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i17  (.D(recv_buffer[30]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[29]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i17 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i16  (.D(recv_buffer[29]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[28]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i16 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i15  (.D(recv_buffer[28]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[27]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i15 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i14  (.D(recv_buffer[27]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[26]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i14 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i13  (.D(recv_buffer[26]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[25]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i13 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i12  (.D(recv_buffer[25]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[24]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i12 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i11  (.D(recv_buffer[24]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[23]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i11 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i10  (.D(recv_buffer[23]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[22]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i10 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i9  (.D(recv_buffer[22]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[21]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i9 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i8  (.D(recv_buffer[21]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[20]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i8 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i7  (.D(recv_buffer[20]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[19]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i7 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i6  (.D(recv_buffer[19]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[18]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i6 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i5  (.D(recv_buffer[18]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[17]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i5 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i4  (.D(recv_buffer[17]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[16]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i4 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i3  (.D(recv_buffer[16]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[15]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i3 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i2  (.D(recv_buffer[15]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[14]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i2 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i1  (.D(recv_buffer[14]), .SP(clkout_c_enable_99), 
            .CK(clkout_c), .Q(recv_buffer[13]));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i1 .GSR = "DISABLED";
    LUT4 i2893_3_lut_4_lut_4_lut (.A(MISOb), .B(n21864), .C(n21865), .D(send_buffer[1]), 
         .Z(MISOb_N_660)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam i2893_3_lut_4_lut_4_lut.init = 16'hf2c2;
    LUT4 mux_51_i53_3_lut_4_lut (.A(send_buffer[53]), .B(n21864), .C(n21865), 
         .D(MISOb_N_666[52]), .Z(send_buffer_95__N_346[52])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i53_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_51_i54_3_lut_4_lut (.A(send_buffer[53]), .B(n21864), .C(n21865), 
         .D(MISOb_N_666[54]), .Z(send_buffer_95__N_346[53])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i54_3_lut_4_lut.init = 16'hf202;
    LUT4 mux_51_i32_3_lut_4_lut (.A(send_buffer[32]), .B(n21864), .C(n21865), 
         .D(MISOb_N_666[31]), .Z(send_buffer_95__N_346[31])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i32_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_51_i33_3_lut_4_lut (.A(send_buffer[32]), .B(n21864), .C(n21865), 
         .D(MISOb_N_666[33]), .Z(send_buffer_95__N_346[32])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i33_3_lut_4_lut.init = 16'hf202;
    LUT4 CSold_I_0_132_2_lut (.A(CSold), .B(CSlatched), .Z(enable_m1_N_633)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(139[7:42])
    defparam CSold_I_0_132_2_lut.init = 16'h8888;
    FD1P3JX speed_set_m3_i0_i5 (.D(recv_buffer[38]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i6 (.D(recv_buffer[39]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i7 (.D(recv_buffer[40]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i8 (.D(recv_buffer[41]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i9 (.D(recv_buffer[42]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i9.GSR = "DISABLED";
    LUT4 mux_51_i8_3_lut_4_lut (.A(send_buffer[7]), .B(n21864), .C(n21865), 
         .D(MISOb_N_666[8]), .Z(send_buffer_95__N_346[7])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i8_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_51_i7_3_lut_4_lut_4_lut (.A(send_buffer[6]), .B(n21864), .C(n21865), 
         .D(send_buffer[7]), .Z(send_buffer_95__N_346[6])) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i7_3_lut_4_lut_4_lut.init = 16'hf2c2;
    LUT4 mux_51_i6_3_lut_4_lut_4_lut (.A(send_buffer[5]), .B(n21864), .C(n21865), 
         .D(send_buffer[6]), .Z(send_buffer_95__N_346[5])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i6_3_lut_4_lut_4_lut.init = 16'h3e0e;
    LUT4 i2_4_lut (.A(n3480), .B(n3456), .C(n39), .D(n40), .Z(enable_m4_N_649)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 mux_51_i5_3_lut_4_lut_4_lut (.A(send_buffer[4]), .B(n21864), .C(n21865), 
         .D(send_buffer[5]), .Z(send_buffer_95__N_346[4])) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i5_3_lut_4_lut_4_lut.init = 16'hf2c2;
    LUT4 mux_51_i4_3_lut_4_lut_4_lut (.A(send_buffer[3]), .B(n21864), .C(n21865), 
         .D(send_buffer[4]), .Z(send_buffer_95__N_346[3])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i4_3_lut_4_lut_4_lut.init = 16'h3e0e;
    LUT4 mux_51_i2_3_lut_4_lut_4_lut (.A(send_buffer[2]), .B(n21864), .C(n21865), 
         .D(send_buffer[1]), .Z(send_buffer_95__N_346[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A (B (C)+!B (C+!(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i2_3_lut_4_lut_4_lut.init = 16'h2f2c;
    LUT4 mux_51_i3_3_lut_4_lut_4_lut (.A(send_buffer[2]), .B(n21864), .C(n21865), 
         .D(send_buffer[3]), .Z(send_buffer_95__N_346[2])) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i3_3_lut_4_lut_4_lut.init = 16'hf2c2;
    LUT4 i18_4_lut (.A(recv_buffer[25]), .B(n36), .C(n28), .D(recv_buffer[24]), 
         .Z(n39)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(recv_buffer[27]), .B(n38), .C(n32), .D(recv_buffer[22]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(n169[0]), .B(recv_buffer[19]), .C(recv_buffer[29]), 
         .D(recv_buffer[23]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(recv_buffer[13]), .B(recv_buffer[14]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i1_4_lut (.A(hallsense_m1[2]), .B(n21919), .C(dir_m1), .D(hallsense_m1[1]), 
         .Z(n2786)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut.init = 16'h4008;
    LUT4 i1_4_lut_adj_132 (.A(hallsense_m1[1]), .B(n21919), .C(dir_m1), 
         .D(hallsense_m1[0]), .Z(n2822)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_132.init = 16'h4008;
    LUT4 i17_4_lut (.A(recv_buffer[20]), .B(n34), .C(n24), .D(recv_buffer[28]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(recv_buffer[18]), .B(recv_buffer[15]), .C(recv_buffer[26]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(recv_buffer[32]), .B(recv_buffer[31]), .C(recv_buffer[21]), 
         .D(recv_buffer[16]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(recv_buffer[30]), .B(recv_buffer[17]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i2_4_lut_adj_133 (.A(n3432), .B(n3408), .C(n39_adj_1874), .D(n40_adj_1875), 
         .Z(enable_m3_N_642)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_133.init = 16'h8880;
    LUT4 i18_4_lut_adj_134 (.A(recv_buffer[46]), .B(n36_adj_1876), .C(n28_adj_1877), 
         .D(recv_buffer[45]), .Z(n39_adj_1874)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_134.init = 16'hfffe;
    LUT4 i19_4_lut_adj_135 (.A(recv_buffer[48]), .B(n38_adj_1878), .C(n32_adj_1879), 
         .D(recv_buffer[43]), .Z(n40_adj_1875)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_135.init = 16'hfffe;
    LUT4 mux_51_i74_3_lut_4_lut (.A(send_buffer[74]), .B(n21864), .C(n21865), 
         .D(MISOb_N_666[73]), .Z(send_buffer_95__N_346[73])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i74_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_51_i75_3_lut_4_lut (.A(send_buffer[74]), .B(n21864), .C(n21865), 
         .D(MISOb_N_666[75]), .Z(send_buffer_95__N_346[74])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i75_3_lut_4_lut.init = 16'hf202;
    LUT4 i1_4_lut_adj_136 (.A(hallsense_m2[2]), .B(n21912), .C(dir_m2), 
         .D(hallsense_m2[1]), .Z(n2916)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_136.init = 16'h4008;
    LUT4 i1_4_lut_adj_137 (.A(hallsense_m2[1]), .B(n21912), .C(dir_m2), 
         .D(hallsense_m2[0]), .Z(n2952)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_137.init = 16'h4008;
    FD1P3IX speed_set_m3_i0_i10 (.D(recv_buffer[43]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i11 (.D(recv_buffer[44]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i12 (.D(recv_buffer[45]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i12.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i13 (.D(recv_buffer[46]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i13.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i14 (.D(recv_buffer[47]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i15 (.D(recv_buffer[48]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i15.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i16 (.D(recv_buffer[49]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i16.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i17 (.D(recv_buffer[50]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i17.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i18 (.D(recv_buffer[51]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i18.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i19 (.D(recv_buffer[52]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i20 (.D(recv_buffer[53]), .SP(clkout_c_enable_245), 
            .CD(n13012), .CK(clkout_c), .Q(speed_set_m3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i20.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i1 (.D(recv_buffer[13]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i1.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i2 (.D(recv_buffer[14]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i2.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i3 (.D(recv_buffer[15]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i4 (.D(recv_buffer[16]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i4.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i5 (.D(recv_buffer[17]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i6 (.D(recv_buffer[18]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i7 (.D(recv_buffer[19]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i8 (.D(recv_buffer[20]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i8.GSR = "DISABLED";
    LUT4 i15_4_lut_adj_138 (.A(recv_buffer[33]), .B(recv_buffer[40]), .C(recv_buffer[50]), 
         .D(recv_buffer[44]), .Z(n36_adj_1876)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_138.init = 16'hfffe;
    LUT4 i7_2_lut_adj_139 (.A(recv_buffer[34]), .B(recv_buffer[35]), .Z(n28_adj_1877)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_139.init = 16'heeee;
    LUT4 i17_4_lut_adj_140 (.A(recv_buffer[41]), .B(n34_adj_1880), .C(n24_adj_1881), 
         .D(recv_buffer[49]), .Z(n38_adj_1878)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_140.init = 16'hfffe;
    LUT4 i11_3_lut_adj_141 (.A(recv_buffer[39]), .B(recv_buffer[36]), .C(recv_buffer[47]), 
         .Z(n32_adj_1879)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_141.init = 16'hfefe;
    LUT4 i13_4_lut_adj_142 (.A(recv_buffer[53]), .B(recv_buffer[52]), .C(recv_buffer[42]), 
         .D(recv_buffer[37]), .Z(n34_adj_1880)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_142.init = 16'hfffe;
    LUT4 i3_2_lut_adj_143 (.A(recv_buffer[51]), .B(recv_buffer[38]), .Z(n24_adj_1881)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_143.init = 16'heeee;
    LUT4 i1_4_lut_adj_144 (.A(hallsense_m3[2]), .B(n21907), .C(dir_m3), 
         .D(hallsense_m3[1]), .Z(n3046)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_144.init = 16'h4008;
    LUT4 i1_4_lut_adj_145 (.A(hallsense_m3[1]), .B(n21907), .C(dir_m3), 
         .D(hallsense_m3[0]), .Z(n3082)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_145.init = 16'h4008;
    FD1P3JX speed_set_m4_i0_i9 (.D(recv_buffer[21]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i9.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i10 (.D(recv_buffer[22]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i11 (.D(recv_buffer[23]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i12 (.D(recv_buffer[24]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i12.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i13 (.D(recv_buffer[25]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i13.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i14 (.D(recv_buffer[26]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i15 (.D(recv_buffer[27]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i15.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i16 (.D(recv_buffer[28]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i16.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i17 (.D(recv_buffer[29]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i17.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i18 (.D(recv_buffer[30]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i18.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i19 (.D(recv_buffer[31]), .SP(clkout_c_enable_245), 
            .PD(n12992), .CK(clkout_c), .Q(speed_set_m4[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i20 (.D(recv_buffer[32]), .SP(clkout_c_enable_245), 
            .CD(n12992), .CK(clkout_c), .Q(speed_set_m4[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i20.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i0 (.D(n169[0]), .SP(clkout_c_enable_245), .PD(n12992), 
            .CK(clkout_c), .Q(speed_set_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i0.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i0 (.D(recv_buffer[33]), .SP(clkout_c_enable_245), 
            .PD(n13012), .CK(clkout_c), .Q(speed_set_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i0.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i0 (.D(recv_buffer[54]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i0.GSR = "DISABLED";
    LUT4 i3_4_lut_rep_515 (.A(SCKold), .B(n22383), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_64)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut_rep_515.init = 16'h0400;
    FD1P3AX send_buffer_i0_i1 (.D(send_buffer_95__N_346[1]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i1.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i2 (.D(send_buffer_95__N_346[2]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i3 (.D(send_buffer_95__N_346[3]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i4 (.D(send_buffer_95__N_346[4]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i4.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i5 (.D(send_buffer_95__N_346[5]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i5.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i6 (.D(send_buffer_95__N_346[6]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i7 (.D(send_buffer_95__N_346[7]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i8 (.D(send_buffer_95__N_346[8]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i8.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i9 (.D(send_buffer_95__N_346[9]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i9.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i10 (.D(send_buffer_95__N_346[10]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i10.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i11 (.D(send_buffer_95__N_346[11]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i11.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i12 (.D(send_buffer_95__N_346[12]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i12.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i13 (.D(send_buffer_95__N_346[13]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i13.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i14 (.D(send_buffer_95__N_346[14]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i14.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i15 (.D(send_buffer_95__N_346[15]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i15.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i16 (.D(send_buffer_95__N_346[16]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i16.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i17 (.D(send_buffer_95__N_346[17]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i17.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i18 (.D(send_buffer_95__N_346[18]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i18.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i19 (.D(send_buffer_95__N_346[19]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i19.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i20 (.D(send_buffer_95__N_346[20]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i20.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i21 (.D(send_buffer_95__N_346[21]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i21.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i22 (.D(send_buffer_95__N_346[22]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i22.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i23 (.D(send_buffer_95__N_346[23]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i23.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i24 (.D(send_buffer_95__N_346[24]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i24.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i25 (.D(send_buffer_95__N_346[25]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i25.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i26 (.D(send_buffer_95__N_346[26]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i26.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i27 (.D(send_buffer_95__N_346[27]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i27.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i28 (.D(send_buffer_95__N_346[28]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i28.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i29 (.D(send_buffer_95__N_346[29]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i29.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i30 (.D(send_buffer_95__N_346[30]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i30.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i31 (.D(send_buffer_95__N_346[31]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i31.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i32 (.D(send_buffer_95__N_346[32]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i32.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i33 (.D(send_buffer_95__N_346[33]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i33.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i34 (.D(send_buffer_95__N_346[34]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i34.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i35 (.D(send_buffer_95__N_346[35]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i35.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i36 (.D(send_buffer_95__N_346[36]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i36.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i37 (.D(send_buffer_95__N_346[37]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i37.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i38 (.D(send_buffer_95__N_346[38]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i38.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i39 (.D(send_buffer_95__N_346[39]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i39.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i40 (.D(send_buffer_95__N_346[40]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i40.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i41 (.D(send_buffer_95__N_346[41]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i41.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i42 (.D(send_buffer_95__N_346[42]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i42.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i43 (.D(send_buffer_95__N_346[43]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i43.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i44 (.D(send_buffer_95__N_346[44]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i44.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i45 (.D(send_buffer_95__N_346[45]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i45.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i46 (.D(send_buffer_95__N_346[46]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i46.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i47 (.D(send_buffer_95__N_346[47]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i47.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i48 (.D(send_buffer_95__N_346[48]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i48.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i49 (.D(send_buffer_95__N_346[49]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i49.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i50 (.D(send_buffer_95__N_346[50]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i50.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i51 (.D(send_buffer_95__N_346[51]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i51.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i52 (.D(send_buffer_95__N_346[52]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i52.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i53 (.D(send_buffer_95__N_346[53]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i53.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i54 (.D(send_buffer_95__N_346[54]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i54.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i55 (.D(send_buffer_95__N_346[55]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i55.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i56 (.D(send_buffer_95__N_346[56]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i56.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i57 (.D(send_buffer_95__N_346[57]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i57.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i58 (.D(send_buffer_95__N_346[58]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i58.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i59 (.D(send_buffer_95__N_346[59]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i59.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i60 (.D(send_buffer_95__N_346[60]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i60.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i61 (.D(send_buffer_95__N_346[61]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i61.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i62 (.D(send_buffer_95__N_346[62]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i62.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i63 (.D(send_buffer_95__N_346[63]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i63.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i64 (.D(send_buffer_95__N_346[64]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i64.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i65 (.D(send_buffer_95__N_346[65]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i65.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i66 (.D(send_buffer_95__N_346[66]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i66.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i67 (.D(send_buffer_95__N_346[67]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i67.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i68 (.D(send_buffer_95__N_346[68]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i68.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i69 (.D(send_buffer_95__N_346[69]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i69.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i70 (.D(send_buffer_95__N_346[70]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i70.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i71 (.D(send_buffer_95__N_346[71]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i71.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i72 (.D(send_buffer_95__N_346[72]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i72.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i73 (.D(send_buffer_95__N_346[73]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i73.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i74 (.D(send_buffer_95__N_346[74]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i74.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i75 (.D(send_buffer_95__N_346[75]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i75.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i76 (.D(send_buffer_95__N_346[76]), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(send_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i76.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i77 (.D(send_buffer_95__N_346[77]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i77.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i78 (.D(send_buffer_95__N_346[78]), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(send_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i78.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i79 (.D(send_buffer_95__N_346[79]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i79.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i80 (.D(send_buffer_95__N_346[80]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i80.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i81 (.D(send_buffer_95__N_346[81]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i81.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i82 (.D(send_buffer_95__N_346[82]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i82.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i83 (.D(send_buffer_95__N_346[83]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i83.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i84 (.D(send_buffer_95__N_346[84]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i84.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i85 (.D(send_buffer_95__N_346[85]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i85.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i86 (.D(send_buffer_95__N_346[86]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i86.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i87 (.D(send_buffer_95__N_346[87]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i87.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i88 (.D(send_buffer_95__N_346[88]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i88.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i89 (.D(send_buffer_95__N_346[89]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i89.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i90 (.D(send_buffer_95__N_346[90]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i90.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i91 (.D(send_buffer_95__N_346[91]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i91.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i92 (.D(send_buffer_95__N_346[92]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i92.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i93 (.D(send_buffer_95__N_346[93]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i93.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i94 (.D(\send_buffer_95__N_346[94] ), .SP(rst), 
            .CK(clkout_c), .Q(\send_buffer[94] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i94.GSR = "DISABLED";
    LUT4 i3_4_lut (.A(SCKold), .B(n22383), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_99)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i1_4_lut_adj_146 (.A(hallsense_m4[2]), .B(n21901), .C(dir_m4), 
         .D(hallsense_m4[1]), .Z(n3176)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_146.init = 16'h4008;
    LUT4 i1_4_lut_adj_147 (.A(hallsense_m4[1]), .B(n21901), .C(dir_m4), 
         .D(hallsense_m4[0]), .Z(n3212)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_147.init = 16'h4008;
    LUT4 MISOb_N_667_bdd_2_lut (.A(MISO_N_624), .B(MISO_N_625), .Z(n21813)) /* synthesis lut_function=(A (B)) */ ;
    defparam MISOb_N_667_bdd_2_lut.init = 16'h8888;
    CCU2D add_16129_16 (.A0(recv_buffer[95]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18895), .S1(n3336));
    defparam add_16129_16.INIT0 = 16'h0aaa;
    defparam add_16129_16.INIT1 = 16'h0000;
    defparam add_16129_16.INJECT1_0 = "NO";
    defparam add_16129_16.INJECT1_1 = "NO";
    CCU2D add_16129_14 (.A0(recv_buffer[93]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[94]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18894), .COUT(n18895));
    defparam add_16129_14.INIT0 = 16'h5aaa;
    defparam add_16129_14.INIT1 = 16'h5aaa;
    defparam add_16129_14.INJECT1_0 = "NO";
    defparam add_16129_14.INJECT1_1 = "NO";
    CCU2D add_16129_12 (.A0(recv_buffer[91]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[92]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18893), .COUT(n18894));
    defparam add_16129_12.INIT0 = 16'h5aaa;
    defparam add_16129_12.INIT1 = 16'h5aaa;
    defparam add_16129_12.INJECT1_0 = "NO";
    defparam add_16129_12.INJECT1_1 = "NO";
    CCU2D add_16129_10 (.A0(recv_buffer[89]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[90]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18892), .COUT(n18893));
    defparam add_16129_10.INIT0 = 16'h5555;
    defparam add_16129_10.INIT1 = 16'h5aaa;
    defparam add_16129_10.INJECT1_0 = "NO";
    defparam add_16129_10.INJECT1_1 = "NO";
    LUT4 SCKold_I_0_2_lut_rep_467 (.A(SCKold), .B(SCKlatched), .Z(n21887)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(193[8:45])
    defparam SCKold_I_0_2_lut_rep_467.init = 16'h2222;
    CCU2D add_16129_8 (.A0(recv_buffer[87]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[88]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18891), .COUT(n18892));
    defparam add_16129_8.INIT0 = 16'h5aaa;
    defparam add_16129_8.INIT1 = 16'h5aaa;
    defparam add_16129_8.INJECT1_0 = "NO";
    defparam add_16129_8.INJECT1_1 = "NO";
    CCU2D add_16129_6 (.A0(recv_buffer[85]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[86]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18890), .COUT(n18891));
    defparam add_16129_6.INIT0 = 16'h5555;
    defparam add_16129_6.INIT1 = 16'h5555;
    defparam add_16129_6.INJECT1_0 = "NO";
    defparam add_16129_6.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_148 (.A(n3336), .B(n3312), .C(n39_adj_1882), .D(n40_adj_1883), 
         .Z(enable_m1_N_627)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_148.init = 16'h8880;
    CCU2D add_16129_4 (.A0(recv_buffer[83]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[84]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18889), .COUT(n18890));
    defparam add_16129_4.INIT0 = 16'h5aaa;
    defparam add_16129_4.INIT1 = 16'h5555;
    defparam add_16129_4.INJECT1_0 = "NO";
    defparam add_16129_4.INJECT1_1 = "NO";
    LUT4 i18_4_lut_adj_149 (.A(recv_buffer[88]), .B(n36_adj_1884), .C(n28_adj_1885), 
         .D(recv_buffer[87]), .Z(n39_adj_1882)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i18_4_lut_adj_149.init = 16'hfffe;
    LUT4 i19_4_lut_adj_150 (.A(recv_buffer[90]), .B(n38_adj_1886), .C(n32_adj_1887), 
         .D(recv_buffer[85]), .Z(n40_adj_1883)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i19_4_lut_adj_150.init = 16'hfffe;
    FD1P3JX speed_set_m1_i0_i1 (.D(recv_buffer[76]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i1.GSR = "DISABLED";
    LUT4 i15_4_lut_adj_151 (.A(recv_buffer[75]), .B(recv_buffer[82]), .C(recv_buffer[92]), 
         .D(recv_buffer[86]), .Z(n36_adj_1884)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i15_4_lut_adj_151.init = 16'hfffe;
    FD1P3JX speed_set_m1_i0_i2 (.D(recv_buffer[77]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i2.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i3 (.D(recv_buffer[78]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i4 (.D(recv_buffer[79]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i4.GSR = "DISABLED";
    LUT4 i7_2_lut_adj_152 (.A(recv_buffer[76]), .B(recv_buffer[77]), .Z(n28_adj_1885)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i7_2_lut_adj_152.init = 16'heeee;
    FD1P3JX speed_set_m1_i0_i5 (.D(recv_buffer[80]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i6 (.D(recv_buffer[81]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i7 (.D(recv_buffer[82]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i8 (.D(recv_buffer[83]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i9 (.D(recv_buffer[84]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i9.GSR = "DISABLED";
    CCU2D add_16129_2 (.A0(recv_buffer[81]), .B0(recv_buffer[80]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[82]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18889));
    defparam add_16129_2.INIT0 = 16'h7000;
    defparam add_16129_2.INIT1 = 16'h5aaa;
    defparam add_16129_2.INJECT1_0 = "NO";
    defparam add_16129_2.INJECT1_1 = "NO";
    FD1P3IX speed_set_m1_i0_i10 (.D(recv_buffer[85]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i11 (.D(recv_buffer[86]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i11.GSR = "DISABLED";
    CCU2D add_16130_21 (.A0(recv_buffer[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18888), .S1(n3408));
    defparam add_16130_21.INIT0 = 16'h5555;
    defparam add_16130_21.INIT1 = 16'h0000;
    defparam add_16130_21.INJECT1_0 = "NO";
    defparam add_16130_21.INJECT1_1 = "NO";
    FD1P3IX speed_set_m1_i0_i12 (.D(recv_buffer[87]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i12.GSR = "DISABLED";
    LUT4 i17_4_lut_adj_153 (.A(recv_buffer[83]), .B(n34_adj_1888), .C(n24_adj_1889), 
         .D(recv_buffer[91]), .Z(n38_adj_1886)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i17_4_lut_adj_153.init = 16'hfffe;
    FD1P3IX speed_set_m1_i0_i13 (.D(recv_buffer[88]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i13.GSR = "DISABLED";
    CCU2D add_16130_19 (.A0(recv_buffer[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18887), .COUT(n18888));
    defparam add_16130_19.INIT0 = 16'hf555;
    defparam add_16130_19.INIT1 = 16'hf555;
    defparam add_16130_19.INJECT1_0 = "NO";
    defparam add_16130_19.INJECT1_1 = "NO";
    FD1P3JX speed_set_m1_i0_i14 (.D(recv_buffer[89]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i14.GSR = "DISABLED";
    LUT4 i11_3_lut_adj_154 (.A(recv_buffer[81]), .B(recv_buffer[78]), .C(recv_buffer[89]), 
         .Z(n32_adj_1887)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i11_3_lut_adj_154.init = 16'hfefe;
    FD1P3IX speed_set_m1_i0_i15 (.D(recv_buffer[90]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i15.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i16 (.D(recv_buffer[91]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i16.GSR = "DISABLED";
    LUT4 i13_4_lut_adj_155 (.A(recv_buffer[95]), .B(recv_buffer[94]), .C(recv_buffer[84]), 
         .D(recv_buffer[79]), .Z(n34_adj_1888)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i13_4_lut_adj_155.init = 16'hfffe;
    LUT4 i3_2_lut_adj_156 (.A(recv_buffer[93]), .B(recv_buffer[80]), .Z(n24_adj_1889)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(146[7:28])
    defparam i3_2_lut_adj_156.init = 16'heeee;
    CCU2D add_16130_17 (.A0(recv_buffer[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18886), .COUT(n18887));
    defparam add_16130_17.INIT0 = 16'hf555;
    defparam add_16130_17.INIT1 = 16'hf555;
    defparam add_16130_17.INJECT1_0 = "NO";
    defparam add_16130_17.INJECT1_1 = "NO";
    CCU2D add_16130_15 (.A0(recv_buffer[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18885), .COUT(n18886));
    defparam add_16130_15.INIT0 = 16'h0aaa;
    defparam add_16130_15.INIT1 = 16'hf555;
    defparam add_16130_15.INJECT1_0 = "NO";
    defparam add_16130_15.INJECT1_1 = "NO";
    CCU2D add_16130_13 (.A0(recv_buffer[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18884), .COUT(n18885));
    defparam add_16130_13.INIT0 = 16'hf555;
    defparam add_16130_13.INIT1 = 16'hf555;
    defparam add_16130_13.INJECT1_0 = "NO";
    defparam add_16130_13.INJECT1_1 = "NO";
    FD1P3AX CSold_113_rep_510 (.D(CSlatched), .SP(clkout_c_enable_219), 
            .CK(clkout_c), .Q(n22382));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_113_rep_510.GSR = "DISABLED";
    CCU2D add_16130_11 (.A0(recv_buffer[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18883), .COUT(n18884));
    defparam add_16130_11.INIT0 = 16'h0aaa;
    defparam add_16130_11.INIT1 = 16'h0aaa;
    defparam add_16130_11.INJECT1_0 = "NO";
    defparam add_16130_11.INJECT1_1 = "NO";
    LUT4 CSlatched_I_0_1_lut_rep_469 (.A(CSlatched), .Z(n21889)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam CSlatched_I_0_1_lut_rep_469.init = 16'h5555;
    CCU2D add_16130_9 (.A0(recv_buffer[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18882), .COUT(n18883));
    defparam add_16130_9.INIT0 = 16'hf555;
    defparam add_16130_9.INIT1 = 16'h0aaa;
    defparam add_16130_9.INJECT1_0 = "NO";
    defparam add_16130_9.INJECT1_1 = "NO";
    LUT4 i13173_3_lut_rep_443_4_lut_4_lut (.A(n22381), .B(\send_buffer[94] ), 
         .C(\speed_m1[19] ), .D(n22382), .Z(n21863)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam i13173_3_lut_rep_443_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_16130_7 (.A0(recv_buffer[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18881), .COUT(n18882));
    defparam add_16130_7.INIT0 = 16'hf555;
    defparam add_16130_7.INIT1 = 16'hf555;
    defparam add_16130_7.INJECT1_0 = "NO";
    defparam add_16130_7.INJECT1_1 = "NO";
    LUT4 CSold_I_0_2_lut_rep_444_2_lut (.A(n22381), .B(n22382), .Z(n21864)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam CSold_I_0_2_lut_rep_444_2_lut.init = 16'h4444;
    CCU2D add_16130_5 (.A0(recv_buffer[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18880), .COUT(n18881));
    defparam add_16130_5.INIT0 = 16'hf555;
    defparam add_16130_5.INIT1 = 16'h0aaa;
    defparam add_16130_5.INJECT1_0 = "NO";
    defparam add_16130_5.INJECT1_1 = "NO";
    LUT4 mux_9_i56_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[55]), .C(\speed_m2[1] ), 
         .D(n22382), .Z(MISOb_N_666[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i57_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[56]), .C(\speed_m2[2] ), 
         .D(n22382), .Z(MISOb_N_666[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3JX speed_set_m1_i0_i17 (.D(recv_buffer[92]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i17.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i18 (.D(recv_buffer[93]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i18.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i19 (.D(recv_buffer[94]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i20 (.D(recv_buffer[95]), .SP(clkout_c_enable_245), 
            .CD(n13052), .CK(clkout_c), .Q(speed_set_m1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i20.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i1 (.D(recv_buffer[55]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i1.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i2 (.D(recv_buffer[56]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i2.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i3 (.D(recv_buffer[57]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i4 (.D(recv_buffer[58]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i4.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i5 (.D(recv_buffer[59]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i6 (.D(recv_buffer[60]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i7 (.D(recv_buffer[61]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i8 (.D(recv_buffer[62]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i9 (.D(recv_buffer[63]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i9.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i10 (.D(recv_buffer[64]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i11 (.D(recv_buffer[65]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i12 (.D(recv_buffer[66]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i12.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i13 (.D(recv_buffer[67]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i13.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i14 (.D(recv_buffer[68]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i15 (.D(recv_buffer[69]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i15.GSR = "DISABLED";
    LUT4 i13185_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[52]), .C(\speed_m3[19] ), 
         .D(n22382), .Z(MISOb_N_666[52])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam i13185_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i58_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[57]), .C(\speed_m2[3] ), 
         .D(n22382), .Z(MISOb_N_666[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i55_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[54]), .C(\speed_m2[0] ), 
         .D(n22382), .Z(MISOb_N_666[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i59_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[58]), .C(\speed_m2[4] ), 
         .D(n22382), .Z(MISOb_N_666[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3JX speed_set_m1_i0_i0 (.D(recv_buffer[75]), .SP(clkout_c_enable_245), 
            .PD(n13052), .CK(clkout_c), .Q(speed_set_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i0.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i16 (.D(recv_buffer[70]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i16.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i17 (.D(recv_buffer[71]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i17.GSR = "DISABLED";
    LUT4 mux_9_i60_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[59]), .C(\speed_m2[5] ), 
         .D(n22382), .Z(MISOb_N_666[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i61_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[60]), .C(\speed_m2[6] ), 
         .D(n22382), .Z(MISOb_N_666[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i62_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[61]), .C(\speed_m2[7] ), 
         .D(n22382), .Z(MISOb_N_666[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_16130_3 (.A0(recv_buffer[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18879), .COUT(n18880));
    defparam add_16130_3.INIT0 = 16'hf555;
    defparam add_16130_3.INIT1 = 16'hf555;
    defparam add_16130_3.INJECT1_0 = "NO";
    defparam add_16130_3.INJECT1_1 = "NO";
    LUT4 mux_9_i63_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[62]), .C(\speed_m2[8] ), 
         .D(n22382), .Z(MISOb_N_666[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i64_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[63]), .C(\speed_m2[9] ), 
         .D(n22382), .Z(MISOb_N_666[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i65_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[64]), .C(\speed_m2[10] ), 
         .D(n22382), .Z(MISOb_N_666[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i66_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[65]), .C(\speed_m2[11] ), 
         .D(n22382), .Z(MISOb_N_666[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i67_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[66]), .C(\speed_m2[12] ), 
         .D(n22382), .Z(MISOb_N_666[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i68_3_lut_4_lut_4_lut (.A(CSlatched), .B(send_buffer[67]), 
         .C(\speed_m2[13] ), .D(CSold), .Z(MISOb_N_666[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i69_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[68]), .C(\speed_m2[14] ), 
         .D(n22382), .Z(MISOb_N_666[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i70_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[69]), .C(\speed_m2[15] ), 
         .D(n22382), .Z(MISOb_N_666[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i71_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[70]), .C(\speed_m2[16] ), 
         .D(n22382), .Z(MISOb_N_666[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i72_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[71]), .C(\speed_m2[17] ), 
         .D(n22382), .Z(MISOb_N_666[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3JX speed_set_m2_i0_i18 (.D(recv_buffer[72]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i18.GSR = "DISABLED";
    CCU2D add_16130_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[33]), .B1(recv_buffer[34]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18879));
    defparam add_16130_1.INIT0 = 16'hF000;
    defparam add_16130_1.INIT1 = 16'ha666;
    defparam add_16130_1.INJECT1_0 = "NO";
    defparam add_16130_1.INJECT1_1 = "NO";
    LUT4 mux_9_i19_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[18]), .C(\speed_m4[6] ), 
         .D(n22382), .Z(MISOb_N_666[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i18_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[17]), .C(\speed_m4[5] ), 
         .D(n22382), .Z(MISOb_N_666[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3JX speed_set_m2_i0_i19 (.D(recv_buffer[73]), .SP(clkout_c_enable_245), 
            .PD(n13032), .CK(clkout_c), .Q(speed_set_m2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i19.GSR = "DISABLED";
    LUT4 mux_9_i73_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[72]), .C(\speed_m2[18] ), 
         .D(n22382), .Z(MISOb_N_666[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i13184_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[73]), .C(\speed_m2[19] ), 
         .D(n22382), .Z(MISOb_N_666[73])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam i13184_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i76_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[75]), .C(\speed_m1[0] ), 
         .D(n22382), .Z(MISOb_N_666[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i77_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[76]), .C(\speed_m1[1] ), 
         .D(n22382), .Z(MISOb_N_666[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i78_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[77]), .C(\speed_m1[2] ), 
         .D(n22382), .Z(MISOb_N_666[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i79_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[78]), .C(\speed_m1[3] ), 
         .D(n22382), .Z(MISOb_N_666[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i80_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[79]), .C(\speed_m1[4] ), 
         .D(n22382), .Z(MISOb_N_666[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i81_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[80]), .C(\speed_m1[5] ), 
         .D(n22382), .Z(MISOb_N_666[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i82_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[81]), .C(\speed_m1[6] ), 
         .D(n22382), .Z(MISOb_N_666[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i83_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[82]), .C(\speed_m1[7] ), 
         .D(n22382), .Z(MISOb_N_666[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i84_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[83]), .C(\speed_m1[8] ), 
         .D(n22382), .Z(MISOb_N_666[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i85_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[84]), .C(\speed_m1[9] ), 
         .D(n22382), .Z(MISOb_N_666[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i86_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[85]), .C(\speed_m1[10] ), 
         .D(n22382), .Z(MISOb_N_666[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i87_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[86]), .C(\speed_m1[11] ), 
         .D(n22382), .Z(MISOb_N_666[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i88_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[87]), .C(\speed_m1[12] ), 
         .D(n22382), .Z(MISOb_N_666[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i89_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[88]), .C(\speed_m1[13] ), 
         .D(n22382), .Z(MISOb_N_666[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i90_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[89]), .C(\speed_m1[14] ), 
         .D(n22382), .Z(MISOb_N_666[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i91_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[90]), .C(\speed_m1[15] ), 
         .D(n22382), .Z(MISOb_N_666[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i92_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[91]), .C(\speed_m1[16] ), 
         .D(n22382), .Z(MISOb_N_666[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i21_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[20]), .C(\speed_m4[8] ), 
         .D(n22382), .Z(MISOb_N_666[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i20_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[19]), .C(\speed_m4[7] ), 
         .D(n22382), .Z(MISOb_N_666[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i93_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[92]), .C(\speed_m1[17] ), 
         .D(n22382), .Z(MISOb_N_666[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i94_3_lut_4_lut_4_lut (.A(CSlatched), .B(send_buffer[93]), 
         .C(\speed_m1[18] ), .D(CSold), .Z(MISOb_N_666[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i23_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[22]), .C(\speed_m4[10] ), 
         .D(n22382), .Z(MISOb_N_666[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i22_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[21]), .C(\speed_m4[9] ), 
         .D(n22382), .Z(MISOb_N_666[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i24_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[23]), .C(\speed_m4[11] ), 
         .D(n22382), .Z(MISOb_N_666[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i25_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[24]), .C(\speed_m4[12] ), 
         .D(n22382), .Z(MISOb_N_666[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i26_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[25]), .C(\speed_m4[13] ), 
         .D(n22382), .Z(MISOb_N_666[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i27_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[26]), .C(\speed_m4[14] ), 
         .D(n22382), .Z(MISOb_N_666[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i28_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[27]), .C(\speed_m4[15] ), 
         .D(n22382), .Z(MISOb_N_666[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i29_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[28]), .C(\speed_m4[16] ), 
         .D(n22382), .Z(MISOb_N_666[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i30_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[29]), .C(\speed_m4[17] ), 
         .D(n22382), .Z(MISOb_N_666[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i31_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[30]), .C(\speed_m4[18] ), 
         .D(n22382), .Z(MISOb_N_666[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i9_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[8]), .C(enable_m4), 
         .D(n22382), .Z(MISOb_N_666[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i13186_3_lut_4_lut_4_lut (.A(CSlatched), .B(send_buffer[31]), .C(\speed_m4[19] ), 
         .D(CSold), .Z(MISOb_N_666[31])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam i13186_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i34_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[33]), .C(\speed_m3[0] ), 
         .D(n22382), .Z(MISOb_N_666[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i35_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[34]), .C(\speed_m3[1] ), 
         .D(n22382), .Z(MISOb_N_666[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i36_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[35]), .C(\speed_m3[2] ), 
         .D(n22382), .Z(MISOb_N_666[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i37_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[36]), .C(\speed_m3[3] ), 
         .D(n22382), .Z(MISOb_N_666[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i38_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[37]), .C(\speed_m3[4] ), 
         .D(n22382), .Z(MISOb_N_666[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i39_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[38]), .C(\speed_m3[5] ), 
         .D(n22382), .Z(MISOb_N_666[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i40_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[39]), .C(\speed_m3[6] ), 
         .D(n22382), .Z(MISOb_N_666[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i41_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[40]), .C(\speed_m3[7] ), 
         .D(n22382), .Z(MISOb_N_666[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i42_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[41]), .C(\speed_m3[8] ), 
         .D(n22382), .Z(MISOb_N_666[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i43_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[42]), .C(\speed_m3[9] ), 
         .D(n22382), .Z(MISOb_N_666[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i2656_1_lut (.A(MISO_N_625), .Z(n4884)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(64[1] 216[13])
    defparam i2656_1_lut.init = 16'h5555;
    LUT4 mux_9_i44_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[43]), .C(\speed_m3[10] ), 
         .D(n22382), .Z(MISOb_N_666[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i45_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[44]), .C(\speed_m3[11] ), 
         .D(n22382), .Z(MISOb_N_666[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i46_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[45]), .C(\speed_m3[12] ), 
         .D(n22382), .Z(MISOb_N_666[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i47_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[46]), .C(\speed_m3[13] ), 
         .D(n22382), .Z(MISOb_N_666[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i48_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[47]), .C(\speed_m3[14] ), 
         .D(n22382), .Z(MISOb_N_666[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i49_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[48]), .C(\speed_m3[15] ), 
         .D(n22382), .Z(MISOb_N_666[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i50_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[49]), .C(\speed_m3[16] ), 
         .D(n22382), .Z(MISOb_N_666[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i51_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[50]), .C(\speed_m3[17] ), 
         .D(n22382), .Z(MISOb_N_666[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i52_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[51]), .C(\speed_m3[18] ), 
         .D(n22382), .Z(MISOb_N_666[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i10_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[9]), .C(enable_m3), 
         .D(n22382), .Z(MISOb_N_666[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i11_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[10]), .C(enable_m2), 
         .D(n22382), .Z(MISOb_N_666[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i12_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[11]), .C(enable_m1), 
         .D(n22382), .Z(MISOb_N_666[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i13_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[12]), .C(\speed_m4[0] ), 
         .D(n22382), .Z(MISOb_N_666[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i14_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[13]), .C(\speed_m4[1] ), 
         .D(n22382), .Z(MISOb_N_666[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i15_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[14]), .C(\speed_m4[2] ), 
         .D(n22382), .Z(MISOb_N_666[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i16_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[15]), .C(\speed_m4[3] ), 
         .D(n22382), .Z(MISOb_N_666[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i17_3_lut_4_lut_4_lut (.A(n22381), .B(send_buffer[16]), .C(\speed_m4[4] ), 
         .D(n22382), .Z(MISOb_N_666[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i68_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[67]), 
         .C(MISOb_N_666[68]), .D(n21887), .Z(send_buffer_95__N_346[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i69_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[68]), 
         .C(MISOb_N_666[69]), .D(n21887), .Z(send_buffer_95__N_346[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i70_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[69]), 
         .C(MISOb_N_666[70]), .D(n21887), .Z(send_buffer_95__N_346[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i71_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[70]), 
         .C(MISOb_N_666[71]), .D(n21887), .Z(send_buffer_95__N_346[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i72_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[71]), 
         .C(MISOb_N_666[72]), .D(n21887), .Z(send_buffer_95__N_346[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i73_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[72]), 
         .C(MISOb_N_666[73]), .D(n21887), .Z(send_buffer_95__N_346[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i76_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[75]), 
         .C(MISOb_N_666[76]), .D(n21887), .Z(send_buffer_95__N_346[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i77_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[76]), 
         .C(MISOb_N_666[77]), .D(n21887), .Z(send_buffer_95__N_346[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i78_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[77]), 
         .C(MISOb_N_666[78]), .D(n21887), .Z(send_buffer_95__N_346[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i79_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[78]), 
         .C(MISOb_N_666[79]), .D(n21887), .Z(send_buffer_95__N_346[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i80_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[79]), 
         .C(MISOb_N_666[80]), .D(n21887), .Z(send_buffer_95__N_346[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i81_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[80]), 
         .C(MISOb_N_666[81]), .D(n21887), .Z(send_buffer_95__N_346[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i82_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[81]), 
         .C(MISOb_N_666[82]), .D(n21887), .Z(send_buffer_95__N_346[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX CSlatched_115_rep_509 (.D(HALL_A_OUT_c_c), .SP(clkout_c_enable_244), 
            .CK(clkout_c), .Q(n22381));   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_115_rep_509.GSR = "DISABLED";
    LUT4 mux_51_i83_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[82]), 
         .C(MISOb_N_666[83]), .D(n21887), .Z(send_buffer_95__N_346[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i84_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[83]), 
         .C(MISOb_N_666[84]), .D(n21887), .Z(send_buffer_95__N_346[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i85_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[84]), 
         .C(MISOb_N_666[85]), .D(n21887), .Z(send_buffer_95__N_346[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i86_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[85]), 
         .C(MISOb_N_666[86]), .D(n21887), .Z(send_buffer_95__N_346[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i87_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[86]), 
         .C(MISOb_N_666[87]), .D(n21887), .Z(send_buffer_95__N_346[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i88_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[87]), 
         .C(MISOb_N_666[88]), .D(n21887), .Z(send_buffer_95__N_346[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i89_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[88]), 
         .C(MISOb_N_666[89]), .D(n21887), .Z(send_buffer_95__N_346[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i90_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[89]), 
         .C(MISOb_N_666[90]), .D(n21887), .Z(send_buffer_95__N_346[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i91_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[90]), 
         .C(MISOb_N_666[91]), .D(n21887), .Z(send_buffer_95__N_346[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i92_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[91]), 
         .C(MISOb_N_666[92]), .D(n21887), .Z(send_buffer_95__N_346[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i93_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[92]), 
         .C(MISOb_N_666[93]), .D(n21887), .Z(send_buffer_95__N_346[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i94_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[93]), 
         .C(n21863), .D(n21887), .Z(send_buffer_95__N_346[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i9_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[8]), 
         .C(MISOb_N_666[9]), .D(n21887), .Z(send_buffer_95__N_346[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i10_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[9]), 
         .C(MISOb_N_666[10]), .D(n21887), .Z(send_buffer_95__N_346[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i11_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[10]), 
         .C(MISOb_N_666[11]), .D(n21887), .Z(send_buffer_95__N_346[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i12_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[11]), 
         .C(MISOb_N_666[12]), .D(n21887), .Z(send_buffer_95__N_346[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i13_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[12]), 
         .C(MISOb_N_666[13]), .D(n21887), .Z(send_buffer_95__N_346[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i14_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[13]), 
         .C(MISOb_N_666[14]), .D(n21887), .Z(send_buffer_95__N_346[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i15_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[14]), 
         .C(MISOb_N_666[15]), .D(n21887), .Z(send_buffer_95__N_346[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i16_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[15]), 
         .C(MISOb_N_666[16]), .D(n21887), .Z(send_buffer_95__N_346[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i17_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[16]), 
         .C(MISOb_N_666[17]), .D(n21887), .Z(send_buffer_95__N_346[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i18_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[17]), 
         .C(MISOb_N_666[18]), .D(n21887), .Z(send_buffer_95__N_346[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i19_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[18]), 
         .C(MISOb_N_666[19]), .D(n21887), .Z(send_buffer_95__N_346[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i20_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[19]), 
         .C(MISOb_N_666[20]), .D(n21887), .Z(send_buffer_95__N_346[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i21_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[20]), 
         .C(MISOb_N_666[21]), .D(n21887), .Z(send_buffer_95__N_346[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i22_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[21]), 
         .C(MISOb_N_666[22]), .D(n21887), .Z(send_buffer_95__N_346[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i23_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[22]), 
         .C(MISOb_N_666[23]), .D(n21887), .Z(send_buffer_95__N_346[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i24_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[23]), 
         .C(MISOb_N_666[24]), .D(n21887), .Z(send_buffer_95__N_346[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i25_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[24]), 
         .C(MISOb_N_666[25]), .D(n21887), .Z(send_buffer_95__N_346[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i26_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[25]), 
         .C(MISOb_N_666[26]), .D(n21887), .Z(send_buffer_95__N_346[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i27_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[26]), 
         .C(MISOb_N_666[27]), .D(n21887), .Z(send_buffer_95__N_346[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i28_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[27]), 
         .C(MISOb_N_666[28]), .D(n21887), .Z(send_buffer_95__N_346[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i29_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[28]), 
         .C(MISOb_N_666[29]), .D(n21887), .Z(send_buffer_95__N_346[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i30_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[29]), 
         .C(MISOb_N_666[30]), .D(n21887), .Z(send_buffer_95__N_346[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i31_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[30]), 
         .C(MISOb_N_666[31]), .D(n21887), .Z(send_buffer_95__N_346[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i34_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[33]), 
         .C(MISOb_N_666[34]), .D(n21887), .Z(send_buffer_95__N_346[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i35_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[34]), 
         .C(MISOb_N_666[35]), .D(n21887), .Z(send_buffer_95__N_346[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i36_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[35]), 
         .C(MISOb_N_666[36]), .D(n21887), .Z(send_buffer_95__N_346[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i37_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[36]), 
         .C(MISOb_N_666[37]), .D(n21887), .Z(send_buffer_95__N_346[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i38_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[37]), 
         .C(MISOb_N_666[38]), .D(n21887), .Z(send_buffer_95__N_346[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i39_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[38]), 
         .C(MISOb_N_666[39]), .D(n21887), .Z(send_buffer_95__N_346[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i40_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[39]), 
         .C(MISOb_N_666[40]), .D(n21887), .Z(send_buffer_95__N_346[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i41_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[40]), 
         .C(MISOb_N_666[41]), .D(n21887), .Z(send_buffer_95__N_346[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i42_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[41]), 
         .C(MISOb_N_666[42]), .D(n21887), .Z(send_buffer_95__N_346[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i43_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[42]), 
         .C(MISOb_N_666[43]), .D(n21887), .Z(send_buffer_95__N_346[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i44_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[43]), 
         .C(MISOb_N_666[44]), .D(n21887), .Z(send_buffer_95__N_346[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i45_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[44]), 
         .C(MISOb_N_666[45]), .D(n21887), .Z(send_buffer_95__N_346[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i46_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[45]), 
         .C(MISOb_N_666[46]), .D(n21887), .Z(send_buffer_95__N_346[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i47_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[46]), 
         .C(MISOb_N_666[47]), .D(n21887), .Z(send_buffer_95__N_346[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i48_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[47]), 
         .C(MISOb_N_666[48]), .D(n21887), .Z(send_buffer_95__N_346[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i49_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[48]), 
         .C(MISOb_N_666[49]), .D(n21887), .Z(send_buffer_95__N_346[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i50_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[49]), 
         .C(MISOb_N_666[50]), .D(n21887), .Z(send_buffer_95__N_346[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i51_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[50]), 
         .C(MISOb_N_666[51]), .D(n21887), .Z(send_buffer_95__N_346[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i52_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[51]), 
         .C(MISOb_N_666[52]), .D(n21887), .Z(send_buffer_95__N_346[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i55_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[54]), 
         .C(MISOb_N_666[55]), .D(n21887), .Z(send_buffer_95__N_346[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i56_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[55]), 
         .C(MISOb_N_666[56]), .D(n21887), .Z(send_buffer_95__N_346[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i57_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[56]), 
         .C(MISOb_N_666[57]), .D(n21887), .Z(send_buffer_95__N_346[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i58_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[57]), 
         .C(MISOb_N_666[58]), .D(n21887), .Z(send_buffer_95__N_346[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i59_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[58]), 
         .C(MISOb_N_666[59]), .D(n21887), .Z(send_buffer_95__N_346[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i60_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[59]), 
         .C(MISOb_N_666[60]), .D(n21887), .Z(send_buffer_95__N_346[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i61_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[60]), 
         .C(MISOb_N_666[61]), .D(n21887), .Z(send_buffer_95__N_346[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i62_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[61]), 
         .C(MISOb_N_666[62]), .D(n21887), .Z(send_buffer_95__N_346[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i63_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[62]), 
         .C(MISOb_N_666[63]), .D(n21887), .Z(send_buffer_95__N_346[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i64_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[63]), 
         .C(MISOb_N_666[64]), .D(n21887), .Z(send_buffer_95__N_346[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i65_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[64]), 
         .C(MISOb_N_666[65]), .D(n21887), .Z(send_buffer_95__N_346[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i66_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[65]), 
         .C(MISOb_N_666[66]), .D(n21887), .Z(send_buffer_95__N_346[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i67_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[66]), 
         .C(MISOb_N_666[67]), .D(n21887), .Z(send_buffer_95__N_346[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i161_2_lut_rep_445_3_lut_3_lut (.A(CSlatched), .B(SCKlatched), 
         .C(SCKold), .Z(n21865)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(117[26:41])
    defparam i161_2_lut_rep_445_3_lut_3_lut.init = 16'h1010;
    CCU2D add_16124_16 (.A0(recv_buffer[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18971), .S1(n3480));
    defparam add_16124_16.INIT0 = 16'h0aaa;
    defparam add_16124_16.INIT1 = 16'h0000;
    defparam add_16124_16.INJECT1_0 = "NO";
    defparam add_16124_16.INJECT1_1 = "NO";
    CCU2D add_16124_14 (.A0(recv_buffer[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18970), .COUT(n18971));
    defparam add_16124_14.INIT0 = 16'h5aaa;
    defparam add_16124_14.INIT1 = 16'h5aaa;
    defparam add_16124_14.INJECT1_0 = "NO";
    defparam add_16124_14.INJECT1_1 = "NO";
    CCU2D add_16124_12 (.A0(recv_buffer[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18969), .COUT(n18970));
    defparam add_16124_12.INIT0 = 16'h5aaa;
    defparam add_16124_12.INIT1 = 16'h5aaa;
    defparam add_16124_12.INJECT1_0 = "NO";
    defparam add_16124_12.INJECT1_1 = "NO";
    CCU2D add_16124_10 (.A0(recv_buffer[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18968), .COUT(n18969));
    defparam add_16124_10.INIT0 = 16'h5555;
    defparam add_16124_10.INIT1 = 16'h5aaa;
    defparam add_16124_10.INJECT1_0 = "NO";
    defparam add_16124_10.INJECT1_1 = "NO";
    CCU2D add_16124_8 (.A0(recv_buffer[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18967), .COUT(n18968));
    defparam add_16124_8.INIT0 = 16'h5aaa;
    defparam add_16124_8.INIT1 = 16'h5aaa;
    defparam add_16124_8.INJECT1_0 = "NO";
    defparam add_16124_8.INJECT1_1 = "NO";
    CCU2D add_16124_6 (.A0(recv_buffer[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18966), .COUT(n18967));
    defparam add_16124_6.INIT0 = 16'h5555;
    defparam add_16124_6.INIT1 = 16'h5555;
    defparam add_16124_6.INJECT1_0 = "NO";
    defparam add_16124_6.INJECT1_1 = "NO";
    CCU2D add_16124_4 (.A0(recv_buffer[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18965), .COUT(n18966));
    defparam add_16124_4.INIT0 = 16'h5aaa;
    defparam add_16124_4.INIT1 = 16'h5555;
    defparam add_16124_4.INJECT1_0 = "NO";
    defparam add_16124_4.INJECT1_1 = "NO";
    CCU2D add_16124_2 (.A0(recv_buffer[18]), .B0(recv_buffer[17]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18965));
    defparam add_16124_2.INIT0 = 16'h7000;
    defparam add_16124_2.INIT1 = 16'h5aaa;
    defparam add_16124_2.INJECT1_0 = "NO";
    defparam add_16124_2.INJECT1_1 = "NO";
    CCU2D add_16125_21 (.A0(recv_buffer[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18964), .S1(n3456));
    defparam add_16125_21.INIT0 = 16'h5555;
    defparam add_16125_21.INIT1 = 16'h0000;
    defparam add_16125_21.INJECT1_0 = "NO";
    defparam add_16125_21.INJECT1_1 = "NO";
    CCU2D add_16125_19 (.A0(recv_buffer[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18963), .COUT(n18964));
    defparam add_16125_19.INIT0 = 16'hf555;
    defparam add_16125_19.INIT1 = 16'hf555;
    defparam add_16125_19.INJECT1_0 = "NO";
    defparam add_16125_19.INJECT1_1 = "NO";
    CCU2D add_16125_17 (.A0(recv_buffer[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18962), .COUT(n18963));
    defparam add_16125_17.INIT0 = 16'hf555;
    defparam add_16125_17.INIT1 = 16'hf555;
    defparam add_16125_17.INJECT1_0 = "NO";
    defparam add_16125_17.INJECT1_1 = "NO";
    CCU2D add_16125_15 (.A0(recv_buffer[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18961), .COUT(n18962));
    defparam add_16125_15.INIT0 = 16'h0aaa;
    defparam add_16125_15.INIT1 = 16'hf555;
    defparam add_16125_15.INJECT1_0 = "NO";
    defparam add_16125_15.INJECT1_1 = "NO";
    CCU2D add_16125_13 (.A0(recv_buffer[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18960), .COUT(n18961));
    defparam add_16125_13.INIT0 = 16'hf555;
    defparam add_16125_13.INIT1 = 16'hf555;
    defparam add_16125_13.INJECT1_0 = "NO";
    defparam add_16125_13.INJECT1_1 = "NO";
    CCU2D add_16125_11 (.A0(recv_buffer[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18959), .COUT(n18960));
    defparam add_16125_11.INIT0 = 16'h0aaa;
    defparam add_16125_11.INIT1 = 16'h0aaa;
    defparam add_16125_11.INJECT1_0 = "NO";
    defparam add_16125_11.INJECT1_1 = "NO";
    CCU2D add_16125_9 (.A0(recv_buffer[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18958), .COUT(n18959));
    defparam add_16125_9.INIT0 = 16'hf555;
    defparam add_16125_9.INIT1 = 16'h0aaa;
    defparam add_16125_9.INJECT1_0 = "NO";
    defparam add_16125_9.INJECT1_1 = "NO";
    CCU2D add_16125_7 (.A0(recv_buffer[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18957), .COUT(n18958));
    defparam add_16125_7.INIT0 = 16'hf555;
    defparam add_16125_7.INIT1 = 16'hf555;
    defparam add_16125_7.INJECT1_0 = "NO";
    defparam add_16125_7.INJECT1_1 = "NO";
    CCU2D add_16125_5 (.A0(recv_buffer[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18956), .COUT(n18957));
    defparam add_16125_5.INIT0 = 16'hf555;
    defparam add_16125_5.INIT1 = 16'h0aaa;
    defparam add_16125_5.INJECT1_0 = "NO";
    defparam add_16125_5.INJECT1_1 = "NO";
    CCU2D add_16125_3 (.A0(recv_buffer[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18955), .COUT(n18956));
    defparam add_16125_3.INIT0 = 16'hf555;
    defparam add_16125_3.INIT1 = 16'hf555;
    defparam add_16125_3.INJECT1_0 = "NO";
    defparam add_16125_3.INJECT1_1 = "NO";
    CCU2D add_16125_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n169[0]), .B1(recv_buffer[13]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18955));
    defparam add_16125_1.INIT0 = 16'hF000;
    defparam add_16125_1.INIT1 = 16'ha666;
    defparam add_16125_1.INJECT1_0 = "NO";
    defparam add_16125_1.INJECT1_1 = "NO";
    CCU2D add_16126_16 (.A0(recv_buffer[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18954), .S1(n3432));
    defparam add_16126_16.INIT0 = 16'h0aaa;
    defparam add_16126_16.INIT1 = 16'h0000;
    defparam add_16126_16.INJECT1_0 = "NO";
    defparam add_16126_16.INJECT1_1 = "NO";
    CCU2D add_16126_14 (.A0(recv_buffer[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18953), .COUT(n18954));
    defparam add_16126_14.INIT0 = 16'h5aaa;
    defparam add_16126_14.INIT1 = 16'h5aaa;
    defparam add_16126_14.INJECT1_0 = "NO";
    defparam add_16126_14.INJECT1_1 = "NO";
    CCU2D add_16126_12 (.A0(recv_buffer[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18952), .COUT(n18953));
    defparam add_16126_12.INIT0 = 16'h5aaa;
    defparam add_16126_12.INIT1 = 16'h5aaa;
    defparam add_16126_12.INJECT1_0 = "NO";
    defparam add_16126_12.INJECT1_1 = "NO";
    CCU2D add_16126_10 (.A0(recv_buffer[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18951), .COUT(n18952));
    defparam add_16126_10.INIT0 = 16'h5555;
    defparam add_16126_10.INIT1 = 16'h5aaa;
    defparam add_16126_10.INJECT1_0 = "NO";
    defparam add_16126_10.INJECT1_1 = "NO";
    CCU2D add_16126_8 (.A0(recv_buffer[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18950), .COUT(n18951));
    defparam add_16126_8.INIT0 = 16'h5aaa;
    defparam add_16126_8.INIT1 = 16'h5aaa;
    defparam add_16126_8.INJECT1_0 = "NO";
    defparam add_16126_8.INJECT1_1 = "NO";
    CCU2D add_16126_6 (.A0(recv_buffer[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18949), .COUT(n18950));
    defparam add_16126_6.INIT0 = 16'h5555;
    defparam add_16126_6.INIT1 = 16'h5555;
    defparam add_16126_6.INJECT1_0 = "NO";
    defparam add_16126_6.INJECT1_1 = "NO";
    CCU2D add_16126_4 (.A0(recv_buffer[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18948), .COUT(n18949));
    defparam add_16126_4.INIT0 = 16'h5aaa;
    defparam add_16126_4.INIT1 = 16'h5555;
    defparam add_16126_4.INJECT1_0 = "NO";
    defparam add_16126_4.INJECT1_1 = "NO";
    CCU2D add_16126_2 (.A0(recv_buffer[39]), .B0(recv_buffer[38]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18948));
    defparam add_16126_2.INIT0 = 16'h7000;
    defparam add_16126_2.INIT1 = 16'h5aaa;
    defparam add_16126_2.INJECT1_0 = "NO";
    defparam add_16126_2.INJECT1_1 = "NO";
    CCU2D add_16118_21 (.A0(recv_buffer[95]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18947), .S1(n3312));
    defparam add_16118_21.INIT0 = 16'h5555;
    defparam add_16118_21.INIT1 = 16'h0000;
    defparam add_16118_21.INJECT1_0 = "NO";
    defparam add_16118_21.INJECT1_1 = "NO";
    CCU2D add_16118_19 (.A0(recv_buffer[93]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[94]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18946), .COUT(n18947));
    defparam add_16118_19.INIT0 = 16'hf555;
    defparam add_16118_19.INIT1 = 16'hf555;
    defparam add_16118_19.INJECT1_0 = "NO";
    defparam add_16118_19.INJECT1_1 = "NO";
    CCU2D add_16118_17 (.A0(recv_buffer[91]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[92]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18945), .COUT(n18946));
    defparam add_16118_17.INIT0 = 16'hf555;
    defparam add_16118_17.INIT1 = 16'hf555;
    defparam add_16118_17.INJECT1_0 = "NO";
    defparam add_16118_17.INJECT1_1 = "NO";
    CCU2D add_16118_15 (.A0(recv_buffer[89]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[90]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18944), .COUT(n18945));
    defparam add_16118_15.INIT0 = 16'h0aaa;
    defparam add_16118_15.INIT1 = 16'hf555;
    defparam add_16118_15.INJECT1_0 = "NO";
    defparam add_16118_15.INJECT1_1 = "NO";
    CCU2D add_16118_13 (.A0(recv_buffer[87]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[88]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18943), .COUT(n18944));
    defparam add_16118_13.INIT0 = 16'hf555;
    defparam add_16118_13.INIT1 = 16'hf555;
    defparam add_16118_13.INJECT1_0 = "NO";
    defparam add_16118_13.INJECT1_1 = "NO";
    CCU2D add_16118_11 (.A0(recv_buffer[85]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[86]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18942), .COUT(n18943));
    defparam add_16118_11.INIT0 = 16'h0aaa;
    defparam add_16118_11.INIT1 = 16'h0aaa;
    defparam add_16118_11.INJECT1_0 = "NO";
    defparam add_16118_11.INJECT1_1 = "NO";
    CCU2D add_16118_9 (.A0(recv_buffer[83]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[84]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18941), .COUT(n18942));
    defparam add_16118_9.INIT0 = 16'hf555;
    defparam add_16118_9.INIT1 = 16'h0aaa;
    defparam add_16118_9.INJECT1_0 = "NO";
    defparam add_16118_9.INJECT1_1 = "NO";
    CCU2D add_16118_7 (.A0(recv_buffer[81]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[82]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18940), .COUT(n18941));
    defparam add_16118_7.INIT0 = 16'hf555;
    defparam add_16118_7.INIT1 = 16'hf555;
    defparam add_16118_7.INJECT1_0 = "NO";
    defparam add_16118_7.INJECT1_1 = "NO";
    CCU2D add_16118_5 (.A0(recv_buffer[79]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[80]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18939), .COUT(n18940));
    defparam add_16118_5.INIT0 = 16'hf555;
    defparam add_16118_5.INIT1 = 16'h0aaa;
    defparam add_16118_5.INJECT1_0 = "NO";
    defparam add_16118_5.INJECT1_1 = "NO";
    CCU2D add_16118_3 (.A0(recv_buffer[77]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[78]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18938), .COUT(n18939));
    defparam add_16118_3.INIT0 = 16'hf555;
    defparam add_16118_3.INIT1 = 16'hf555;
    defparam add_16118_3.INJECT1_0 = "NO";
    defparam add_16118_3.INJECT1_1 = "NO";
    CCU2D add_16118_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[75]), .B1(recv_buffer[76]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18938));
    defparam add_16118_1.INIT0 = 16'hF000;
    defparam add_16118_1.INIT1 = 16'ha666;
    defparam add_16118_1.INJECT1_0 = "NO";
    defparam add_16118_1.INJECT1_1 = "NO";
    CCU2D add_16127_16 (.A0(recv_buffer[74]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18937), .S1(n3384));
    defparam add_16127_16.INIT0 = 16'h0aaa;
    defparam add_16127_16.INIT1 = 16'h0000;
    defparam add_16127_16.INJECT1_0 = "NO";
    defparam add_16127_16.INJECT1_1 = "NO";
    CCU2D add_16127_14 (.A0(recv_buffer[72]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[73]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18936), .COUT(n18937));
    defparam add_16127_14.INIT0 = 16'h5aaa;
    defparam add_16127_14.INIT1 = 16'h5aaa;
    defparam add_16127_14.INJECT1_0 = "NO";
    defparam add_16127_14.INJECT1_1 = "NO";
    CCU2D add_16127_12 (.A0(recv_buffer[70]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[71]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18935), .COUT(n18936));
    defparam add_16127_12.INIT0 = 16'h5aaa;
    defparam add_16127_12.INIT1 = 16'h5aaa;
    defparam add_16127_12.INJECT1_0 = "NO";
    defparam add_16127_12.INJECT1_1 = "NO";
    FD1P3IX speed_set_m2_i0_i20 (.D(recv_buffer[74]), .SP(clkout_c_enable_245), 
            .CD(n13032), .CK(clkout_c), .Q(speed_set_m2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i20.GSR = "DISABLED";
    CCU2D add_16127_10 (.A0(recv_buffer[68]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[69]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18934), .COUT(n18935));
    defparam add_16127_10.INIT0 = 16'h5555;
    defparam add_16127_10.INIT1 = 16'h5aaa;
    defparam add_16127_10.INJECT1_0 = "NO";
    defparam add_16127_10.INJECT1_1 = "NO";
    CCU2D add_16127_8 (.A0(recv_buffer[66]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[67]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18933), .COUT(n18934));
    defparam add_16127_8.INIT0 = 16'h5aaa;
    defparam add_16127_8.INIT1 = 16'h5aaa;
    defparam add_16127_8.INJECT1_0 = "NO";
    defparam add_16127_8.INJECT1_1 = "NO";
    CCU2D add_16127_6 (.A0(recv_buffer[64]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[65]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18932), .COUT(n18933));
    defparam add_16127_6.INIT0 = 16'h5555;
    defparam add_16127_6.INIT1 = 16'h5555;
    defparam add_16127_6.INJECT1_0 = "NO";
    defparam add_16127_6.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_481 (.A(enable_m4), .B(free_m4), .Z(n21901)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_481.init = 16'h2222;
    LUT4 i18371_3_lut_4_lut (.A(enable_m4), .B(free_m4), .C(hallsense_m4[2]), 
         .D(hallsense_m4[0]), .Z(n20030)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i18371_3_lut_4_lut.init = 16'hfddf;
    CCU2D add_16127_4 (.A0(recv_buffer[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18931), .COUT(n18932));
    defparam add_16127_4.INIT0 = 16'h5aaa;
    defparam add_16127_4.INIT1 = 16'h5555;
    defparam add_16127_4.INJECT1_0 = "NO";
    defparam add_16127_4.INJECT1_1 = "NO";
    CCU2D add_16127_2 (.A0(recv_buffer[60]), .B0(recv_buffer[59]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18931));
    defparam add_16127_2.INIT0 = 16'h7000;
    defparam add_16127_2.INIT1 = 16'h5aaa;
    defparam add_16127_2.INJECT1_0 = "NO";
    defparam add_16127_2.INJECT1_1 = "NO";
    CCU2D add_16128_21 (.A0(recv_buffer[74]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18930), .S1(n3360));
    defparam add_16128_21.INIT0 = 16'h5555;
    defparam add_16128_21.INIT1 = 16'h0000;
    defparam add_16128_21.INJECT1_0 = "NO";
    defparam add_16128_21.INJECT1_1 = "NO";
    CCU2D add_16128_19 (.A0(recv_buffer[72]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[73]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18929), .COUT(n18930));
    defparam add_16128_19.INIT0 = 16'hf555;
    defparam add_16128_19.INIT1 = 16'hf555;
    defparam add_16128_19.INJECT1_0 = "NO";
    defparam add_16128_19.INJECT1_1 = "NO";
    CCU2D add_16128_17 (.A0(recv_buffer[70]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[71]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18928), .COUT(n18929));
    defparam add_16128_17.INIT0 = 16'hf555;
    defparam add_16128_17.INIT1 = 16'hf555;
    defparam add_16128_17.INJECT1_0 = "NO";
    defparam add_16128_17.INJECT1_1 = "NO";
    CCU2D add_16128_15 (.A0(recv_buffer[68]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[69]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18927), .COUT(n18928));
    defparam add_16128_15.INIT0 = 16'h0aaa;
    defparam add_16128_15.INIT1 = 16'hf555;
    defparam add_16128_15.INJECT1_0 = "NO";
    defparam add_16128_15.INJECT1_1 = "NO";
    CCU2D add_16128_13 (.A0(recv_buffer[66]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[67]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18926), .COUT(n18927));
    defparam add_16128_13.INIT0 = 16'hf555;
    defparam add_16128_13.INIT1 = 16'hf555;
    defparam add_16128_13.INJECT1_0 = "NO";
    defparam add_16128_13.INJECT1_1 = "NO";
    CCU2D add_16128_11 (.A0(recv_buffer[64]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[65]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18925), .COUT(n18926));
    defparam add_16128_11.INIT0 = 16'h0aaa;
    defparam add_16128_11.INIT1 = 16'h0aaa;
    defparam add_16128_11.INJECT1_0 = "NO";
    defparam add_16128_11.INJECT1_1 = "NO";
    CCU2D add_16128_9 (.A0(recv_buffer[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18924), .COUT(n18925));
    defparam add_16128_9.INIT0 = 16'hf555;
    defparam add_16128_9.INIT1 = 16'h0aaa;
    defparam add_16128_9.INJECT1_0 = "NO";
    defparam add_16128_9.INJECT1_1 = "NO";
    CCU2D add_16128_7 (.A0(recv_buffer[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18923), .COUT(n18924));
    defparam add_16128_7.INIT0 = 16'hf555;
    defparam add_16128_7.INIT1 = 16'hf555;
    defparam add_16128_7.INJECT1_0 = "NO";
    defparam add_16128_7.INJECT1_1 = "NO";
    CCU2D add_16128_5 (.A0(recv_buffer[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18922), .COUT(n18923));
    defparam add_16128_5.INIT0 = 16'hf555;
    defparam add_16128_5.INIT1 = 16'h0aaa;
    defparam add_16128_5.INJECT1_0 = "NO";
    defparam add_16128_5.INJECT1_1 = "NO";
    CCU2D add_16128_3 (.A0(recv_buffer[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18921), .COUT(n18922));
    defparam add_16128_3.INIT0 = 16'hf555;
    defparam add_16128_3.INIT1 = 16'hf555;
    defparam add_16128_3.INJECT1_0 = "NO";
    defparam add_16128_3.INJECT1_1 = "NO";
    CCU2D add_16128_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[54]), .B1(recv_buffer[55]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18921));
    defparam add_16128_1.INIT0 = 16'hF000;
    defparam add_16128_1.INIT1 = 16'ha666;
    defparam add_16128_1.INJECT1_0 = "NO";
    defparam add_16128_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_492 (.A(enable_m2), .B(free_m2), .Z(n21912)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_492.init = 16'h2222;
    PFUMX i18448 (.BLUT(n21813), .ALUT(n21812), .C0(n22383), .Z(MISO_N_670));
    LUT4 i18345_3_lut_4_lut (.A(enable_m2), .B(free_m2), .C(hallsense_m2[2]), 
         .D(hallsense_m2[0]), .Z(n20041)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i18345_3_lut_4_lut.init = 16'hfddf;
    LUT4 i2_3_lut_rep_494 (.A(CSlatched), .B(CSold), .C(n22383), .Z(clkout_c_enable_245)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(139[7:42])
    defparam i2_3_lut_rep_494.init = 16'h8080;
    LUT4 i10765_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22383), .D(enable_m1_N_627), 
         .Z(n13052)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(139[7:42])
    defparam i10765_2_lut_4_lut.init = 16'h0080;
    LUT4 i10745_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22383), .D(enable_m2_N_635), 
         .Z(n13032)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(139[7:42])
    defparam i10745_2_lut_4_lut.init = 16'h0080;
    LUT4 i10705_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22383), .D(enable_m4_N_649), 
         .Z(n12992)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(139[7:42])
    defparam i10705_2_lut_4_lut.init = 16'h0080;
    LUT4 i2_4_lut_adj_157 (.A(n3384), .B(n3360), .C(n39_adj_1898), .D(n40_adj_1899), 
         .Z(enable_m2_N_635)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_157.init = 16'h8880;
    LUT4 i10725_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22383), .D(enable_m3_N_642), 
         .Z(n13012)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/spi loopbacktest v2.vhd(139[7:42])
    defparam i10725_2_lut_4_lut.init = 16'h0080;
    LUT4 i18_4_lut_adj_158 (.A(recv_buffer[67]), .B(n36_adj_1900), .C(n28_adj_1901), 
         .D(recv_buffer[66]), .Z(n39_adj_1898)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_158.init = 16'hfffe;
    LUT4 i19_4_lut_adj_159 (.A(recv_buffer[69]), .B(n38_adj_1902), .C(n32_adj_1903), 
         .D(recv_buffer[64]), .Z(n40_adj_1899)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_159.init = 16'hfffe;
    LUT4 i15_4_lut_adj_160 (.A(recv_buffer[54]), .B(recv_buffer[61]), .C(recv_buffer[71]), 
         .D(recv_buffer[65]), .Z(n36_adj_1900)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_160.init = 16'hfffe;
    LUT4 i7_2_lut_adj_161 (.A(recv_buffer[55]), .B(recv_buffer[56]), .Z(n28_adj_1901)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_161.init = 16'heeee;
    LUT4 i17_4_lut_adj_162 (.A(recv_buffer[62]), .B(n34_adj_1904), .C(n24_adj_1905), 
         .D(recv_buffer[70]), .Z(n38_adj_1902)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_162.init = 16'hfffe;
    LUT4 i3_2_lut_adj_163 (.A(recv_buffer[72]), .B(recv_buffer[59]), .Z(n24_adj_1905)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_163.init = 16'heeee;
    LUT4 i13_4_lut_adj_164 (.A(recv_buffer[74]), .B(recv_buffer[73]), .C(recv_buffer[63]), 
         .D(recv_buffer[58]), .Z(n34_adj_1904)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_164.init = 16'hfffe;
    LUT4 i11_3_lut_adj_165 (.A(recv_buffer[60]), .B(recv_buffer[57]), .C(recv_buffer[68]), 
         .Z(n32_adj_1903)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_165.init = 16'hfefe;
    
endmodule
//
// Verilog Description of module HALL
//

module HALL (clk_1mhz, \speed_m4[0] , clkout_c_enable_244, hallsense_m4, 
            H_A_m4_c, H_B_m4_c, H_C_m4_c, clkout_c_enable_219, GND_net, 
            \speed_m4[1] , \speed_m4[2] , \speed_m4[3] , \speed_m4[4] , 
            \speed_m4[5] , \speed_m4[6] , \speed_m4[7] , \speed_m4[8] , 
            \speed_m4[9] , \speed_m4[10] , \speed_m4[11] , \speed_m4[12] , 
            \speed_m4[13] , \speed_m4[14] , \speed_m4[15] , \speed_m4[16] , 
            \speed_m4[17] , \speed_m4[18] , \speed_m4[19] , n22378);
    input clk_1mhz;
    output \speed_m4[0] ;
    input clkout_c_enable_244;
    output [2:0]hallsense_m4;
    input H_A_m4_c;
    input H_B_m4_c;
    input H_C_m4_c;
    input clkout_c_enable_219;
    input GND_net;
    output \speed_m4[1] ;
    output \speed_m4[2] ;
    output \speed_m4[3] ;
    output \speed_m4[4] ;
    output \speed_m4[5] ;
    output \speed_m4[6] ;
    output \speed_m4[7] ;
    output \speed_m4[8] ;
    output \speed_m4[9] ;
    output \speed_m4[10] ;
    output \speed_m4[11] ;
    output \speed_m4[12] ;
    output \speed_m4[13] ;
    output \speed_m4[14] ;
    output \speed_m4[15] ;
    output \speed_m4[16] ;
    output \speed_m4[17] ;
    output \speed_m4[18] ;
    output \speed_m4[19] ;
    input n22378;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // c:/users/gebruiker/workspace/lattice/final code software/toplevelfinal.vhd(86[9:17])
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_52, n4330;
    wire [19:0]n7;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(62[10:22])
    
    wire stable_counting, n19077;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_old, hall3_lat, hall1_lat, hall2_lat, hall1_old, hall2_old, 
        n21843, n21823, n20082;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(60[10:15])
    
    wire n20305, n21860, n21830, n21825, n20127, n20128, n20129, 
        n20130, n20131, n20132, n20181, n18_adj_1870, n20_adj_1871, 
        n20405, n20263, n20415, n18753, n20377, n18752, n18751, 
        n18750, n18749, n18748, n21879, n21831, n20285;
    wire [6:0]n83;
    
    wire stable_counting_N_1746, n20035, n18_adj_1872, n21916, n15_adj_1873, 
        n18747, n18746, n20361, n18745, n18744, n4, n21915, n21878, 
        n21859;
    
    FD1P3IX speedt__i0 (.D(n7[0]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    FD1P3AX stable_count__i0 (.D(n19077), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m4_c), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m4_c), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m4_c), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_244), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_219), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 i18271_2_lut_rep_402_3_lut_3_lut (.A(n21843), .B(n21823), .C(stable_counting), 
         .Z(clk_1mhz_enable_52)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i18271_2_lut_rep_402_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i1_4_lut_rep_423 (.A(n20082), .B(count[5]), .C(n20305), .D(count[2]), 
         .Z(n21843)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(87[7:21])
    defparam i1_4_lut_rep_423.init = 16'hbfff;
    LUT4 i2497_3_lut_rep_410_4_lut (.A(stable_count[4]), .B(n21860), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n21830)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2497_3_lut_rep_410_4_lut.init = 16'h7f80;
    LUT4 i17449_2_lut_rep_405_4_lut_3_lut_4_lut (.A(stable_count[4]), .B(n21860), 
         .C(stable_count[6]), .D(stable_count[5]), .Z(n21825)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i17449_2_lut_rep_405_4_lut_3_lut_4_lut.init = 16'h7ff8;
    FD1P3AX stable_count__i6 (.D(n20127), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3AX stable_count__i5 (.D(n20128), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3AX stable_count__i4 (.D(n20129), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3AX stable_count__i3 (.D(n20130), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3AX stable_count__i2 (.D(n20131), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3AX stable_count__i1 (.D(n20132), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX speedt__i1 (.D(n7[1]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    FD1P3IX speedt__i2 (.D(n7[2]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n7[3]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n7[4]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n7[5]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n7[6]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n7[7]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n7[8]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n7[9]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n7[10]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n7[11]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n7[12]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n7[13]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n7[14]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n7[15]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n7[16]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n7[17]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n7[18]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n7[19]), .SP(clk_1mhz_enable_52), .CD(n4330), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n7[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    LUT4 i9_4_lut (.A(n20181), .B(n18_adj_1870), .C(count[2]), .D(count[1]), 
         .Z(n20_adj_1871)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i17589_4_lut (.A(count[11]), .B(n20405), .C(n20263), .D(n21825), 
         .Z(n20415)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17589_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(count[5]), .B(count[4]), .C(stable_counting), .D(count[16]), 
         .Z(n18_adj_1870)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18753), 
          .S0(n7[19]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    LUT4 i17579_4_lut (.A(count[12]), .B(n20377), .C(count[0]), .D(count[6]), 
         .Z(n20405)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17579_4_lut.init = 16'hfffe;
    FD1S3IX count__i2 (.D(n7[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n7[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n7[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n7[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n7[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n7[7]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n7[8]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n7[9]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n7[10]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n7[11]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n7[12]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n7[13]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n7[14]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n7[15]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n7[16]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n7[17]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n7[18]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n7[19]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    LUT4 i17439_2_lut (.A(count[8]), .B(count[13]), .Z(n20263)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17439_2_lut.init = 16'heeee;
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18752), .COUT(n18753), .S0(n7[17]), .S1(n7[18]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18751), .COUT(n18752), .S0(n7[15]), .S1(n7[16]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18750), .COUT(n18751), .S0(n7[13]), .S1(n7[14]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18749), .COUT(n18750), .S0(n7[11]), .S1(n7[12]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18748), .COUT(n18749), .S0(n7[9]), .S1(n7[10]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    LUT4 i2490_2_lut_rep_411_3_lut_4_lut (.A(stable_count[3]), .B(n21879), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21831)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2490_2_lut_rep_411_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4_4_lut (.A(n20285), .B(n83[4]), .C(stable_counting_N_1746), 
         .D(stable_count[0]), .Z(n20181)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[7:23])
    defparam i4_4_lut.init = 16'h0100;
    LUT4 mux_28_i2_4_lut (.A(n7[1]), .B(speedt[1]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hac0a;
    LUT4 mux_28_i3_4_lut (.A(n7[2]), .B(speedt[2]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hac0a;
    LUT4 mux_28_i4_4_lut (.A(n7[3]), .B(speedt[3]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hac0a;
    LUT4 i2462_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n83[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2462_2_lut.init = 16'h6666;
    LUT4 mux_28_i5_4_lut (.A(n7[4]), .B(speedt[4]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hac0a;
    LUT4 mux_28_i6_4_lut (.A(n7[5]), .B(speedt[5]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hac0a;
    LUT4 i17481_3_lut (.A(n20035), .B(count[3]), .C(count[17]), .Z(n20305)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17481_3_lut.init = 16'h8080;
    LUT4 mux_28_i7_4_lut (.A(n7[6]), .B(speedt[6]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hac0a;
    LUT4 mux_28_i8_4_lut (.A(n7[7]), .B(speedt[7]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hac0a;
    LUT4 i3_4_lut (.A(count[19]), .B(count[9]), .C(count[14]), .D(count[18]), 
         .Z(n20035)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 mux_28_i9_4_lut (.A(n7[8]), .B(speedt[8]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hac0a;
    LUT4 mux_28_i10_4_lut (.A(n7[9]), .B(speedt[9]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hac0a;
    LUT4 mux_28_i11_4_lut (.A(n7[10]), .B(speedt[10]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hac0a;
    LUT4 mux_28_i12_4_lut (.A(n7[11]), .B(speedt[11]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hac0a;
    LUT4 i9_4_lut_adj_126 (.A(count[0]), .B(n18_adj_1872), .C(n21916), 
         .D(count[12]), .Z(n20082)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(87[7:21])
    defparam i9_4_lut_adj_126.init = 16'hfffe;
    LUT4 i8_4_lut (.A(n15_adj_1873), .B(count[7]), .C(n20263), .D(count[6]), 
         .Z(n18_adj_1872)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(87[7:21])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut (.A(count[11]), .B(count[4]), .C(count[16]), .D(count[1]), 
         .Z(n15_adj_1873)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(87[7:21])
    defparam i5_4_lut.init = 16'hbfff;
    LUT4 mux_28_i13_4_lut (.A(n7[12]), .B(speedt[12]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hac0a;
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    LUT4 mux_28_i14_4_lut (.A(n7[13]), .B(speedt[13]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hac0a;
    LUT4 mux_28_i15_4_lut (.A(n7[14]), .B(speedt[14]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hac0a;
    LUT4 mux_28_i16_4_lut (.A(n7[15]), .B(speedt[15]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hac0a;
    LUT4 mux_28_i17_4_lut (.A(n7[16]), .B(speedt[16]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hac0a;
    LUT4 mux_28_i18_4_lut (.A(n7[17]), .B(speedt[17]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hac0a;
    LUT4 mux_28_i19_4_lut (.A(n7[18]), .B(speedt[18]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hac0a;
    LUT4 mux_28_i20_4_lut (.A(n7[19]), .B(speedt[19]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hac0a;
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18747), 
          .COUT(n18748), .S0(n7[7]), .S1(n7[8]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18746), 
          .COUT(n18747), .S0(n7[5]), .S1(n7[6]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    FD1P3IX stable_counting_62 (.D(n22378), .SP(stable_counting_N_1746), 
            .CD(n20361), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(n7[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_52), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18745), 
          .COUT(n18746), .S0(n7[3]), .S1(n7[4]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18744), 
          .COUT(n18745), .S0(n7[1]), .S1(n7[2]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    LUT4 i2_3_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(92[7:87])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(hall2_old), .B(hall1_old), .C(hall2_lat), .D(hall1_lat), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(92[7:87])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i17536_3_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(n21823), .Z(n20361)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i17536_3_lut.init = 16'hc8c8;
    LUT4 mux_28_i1_4_lut (.A(n7[0]), .B(speedt[0]), .C(n21823), .D(n21843), 
         .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hac0a;
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18744), 
          .S1(n7[0]));   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i2483_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21915), .C(stable_count[4]), 
         .D(stable_count[3]), .Z(n83[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2483_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i10_4_lut_4_lut (.A(clk_1mhz_enable_52), .B(n20415), .C(n20_adj_1871), 
         .D(n20305), .Z(n4330)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i10_4_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_counting), .B(n21823), .C(n21878), 
         .D(stable_counting_N_1746), .Z(n20131)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_127 (.A(stable_counting), .B(n21823), 
         .C(n21859), .D(stable_counting_N_1746), .Z(n20130)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_127.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_128 (.A(stable_counting), .B(n21823), 
         .C(n21830), .D(stable_counting_N_1746), .Z(n20127)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_128.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_129 (.A(stable_counting), .B(n21823), 
         .C(n83[4]), .D(stable_counting_N_1746), .Z(n20129)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_129.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_130 (.A(stable_counting), .B(n21823), 
         .C(n83[1]), .D(stable_counting_N_1746), .Z(n20132)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_130.init = 16'h0070;
    LUT4 i18351_3_lut_4_lut (.A(stable_counting), .B(n21823), .C(stable_counting_N_1746), 
         .D(stable_count[0]), .Z(n19077)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i18351_3_lut_4_lut.init = 16'h0007;
    LUT4 i1_2_lut_3_lut_4_lut_adj_131 (.A(stable_counting), .B(n21823), 
         .C(n21831), .D(stable_counting_N_1746), .Z(n20128)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut_4_lut_adj_131.init = 16'h0070;
    LUT4 i2_3_lut_rep_403_4_lut (.A(n21831), .B(n21830), .C(n83[1]), .D(n20181), 
         .Z(n21823)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_rep_403_4_lut.init = 16'h1000;
    LUT4 i2464_2_lut_rep_495 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21915)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2464_2_lut_rep_495.init = 16'h8888;
    LUT4 i2469_2_lut_rep_458_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21878)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2469_2_lut_rep_458_3_lut.init = 16'h7878;
    LUT4 i2471_2_lut_rep_459_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21879)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2471_2_lut_rep_459_3_lut.init = 16'h8080;
    LUT4 i2478_2_lut_rep_440_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21860)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2478_2_lut_rep_440_3_lut_4_lut.init = 16'h8000;
    LUT4 i2476_2_lut_rep_439_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21859)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i2476_2_lut_rep_439_3_lut_4_lut.init = 16'h78f0;
    LUT4 i17461_2_lut_3_lut_4_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n20285)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/hallinput.vhd(99[21:33])
    defparam i17461_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h7ff8;
    LUT4 i17447_2_lut_rep_496 (.A(count[10]), .B(count[15]), .Z(n21916)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17447_2_lut_rep_496.init = 16'heeee;
    LUT4 i17551_3_lut_4_lut (.A(count[10]), .B(count[15]), .C(stable_count[1]), 
         .D(count[7]), .Z(n20377)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17551_3_lut_4_lut.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module \PID(16000000,160000000,10000000) 
//

module \PID(16000000,160000000,10000000)  (clk_N_683, GND_net, n4201, 
            n4200, intgOut3, backOut2, backOut3, \subOut_24__N_1135[0] , 
            n4203, n4202, dir_m2, dir_m3, dir_m1, dir_m4, n21851, 
            n21835, \speed_m4[3] , n4133, \speed_m4[7] , \speed_m4[8] , 
            \speed_m4[9] , \speed_m4[12] , speed_set_m2, speed_set_m3, 
            n20537, n4204, n10, n10_adj_1, VCC_net, n32, n10_adj_2, 
            n10_adj_3, n10_adj_4, n21, n21_adj_5, n21_adj_6, n21_adj_7, 
            n19454, n21_adj_8, n30, \subOut_24__N_1135[1] , \subOut_24__N_1135[2] , 
            \subOut_24__N_1135[3] , \subOut_24__N_1135[4] , \subOut_24__N_1135[5] , 
            \subOut_24__N_1135[6] , \subOut_24__N_1135[7] , \subOut_24__N_1135[8] , 
            \subOut_24__N_1135[9] , \subOut_24__N_1135[10] , \subOut_24__N_1135[11] , 
            \subOut_24__N_1135[12] , \subOut_24__N_1135[13] , \subOut_24__N_1135[14] , 
            \subOut_24__N_1135[15] , \subOut_24__N_1135[16] , \subOut_24__N_1135[17] , 
            \subOut_24__N_1135[18] , \subOut_24__N_1135[19] , \subOut_24__N_1135[20] , 
            \subOut_24__N_1135[21] , \subOut_24__N_1135[24] , \speed_m1[3] , 
            speed_set_m1, speed_set_m4, \speed_m1[7] , \speed_m1[8] , 
            \speed_m1[9] , \speed_m1[12] , \speed_m1[19] , \speed_m2[19] , 
            n5, \speed_m1[1] , \speed_m2[1] , \speed_m1[2] , \speed_m2[2] , 
            \speed_m1[4] , \speed_m2[4] , \speed_m1[5] , \speed_m2[5] , 
            \speed_m1[6] , \speed_m2[6] , \speed_m1[10] , \speed_m2[10] , 
            \speed_m1[11] , \speed_m2[11] , \speed_m1[13] , \speed_m2[13] , 
            \speed_m1[14] , \speed_m2[14] , \speed_m1[15] , \speed_m2[15] , 
            \speed_m1[16] , \speed_m2[16] , \speed_m1[17] , \speed_m2[17] , 
            \speed_m1[18] , \speed_m2[18] , \speed_m1[0] , \speed_m2[0] , 
            PWMdut_m4, PWMdut_m3, \speed_m3[3] , \speed_m2[3] , n20525, 
            \speed_m3[7] , \speed_m2[7] , \speed_m3[8] , \speed_m2[8] , 
            \speed_m3[9] , \speed_m2[9] , \speed_m3[12] , \speed_m2[12] , 
            \speed_m4[1] , \speed_m3[1] , n21857, \speed_m4[2] , \speed_m3[2] , 
            \speed_m4[4] , \speed_m3[4] , \speed_m4[5] , \speed_m3[5] , 
            \speed_m4[6] , \speed_m3[6] , \speed_m4[10] , \speed_m3[10] , 
            \speed_m4[11] , \speed_m3[11] , \speed_m4[13] , \speed_m3[13] , 
            \speed_m4[14] , \speed_m3[14] , \speed_m4[15] , \speed_m3[15] , 
            \speed_m4[16] , \speed_m3[16] , \speed_m4[17] , \speed_m3[17] , 
            \speed_m4[18] , \speed_m3[18] , \speed_m4[0] , \speed_m3[0] , 
            PWMdut_m2, n9, PWMdut_m1, n20586, n22383, n4208, n7, 
            n4210, n4209, n4212, n4211, n4214, n4213, n4216, n4215, 
            n4218, n4217, n4220, n4219, n4222, n4221, n4224, n4223, 
            n4226, n4225, n4228, n4227, n4229, n4183, n4182, n13, 
            n4185, n4184, n13_adj_9, n13_adj_10, n4187, n4186, n13_adj_11, 
            n13_adj_12, n4189, n4188, n14, n4191, n4190, n4193, 
            n4192, n4195, n4194, n4197, n4196, n4199, n4198);
    input clk_N_683;
    input GND_net;
    output n4201;
    output n4200;
    output [28:0]intgOut3;
    output [28:0]backOut2;
    output [28:0]backOut3;
    input \subOut_24__N_1135[0] ;
    output n4203;
    output n4202;
    output dir_m2;
    output dir_m3;
    output dir_m1;
    output dir_m4;
    output n21851;
    output n21835;
    input \speed_m4[3] ;
    output n4133;
    input \speed_m4[7] ;
    input \speed_m4[8] ;
    input \speed_m4[9] ;
    input \speed_m4[12] ;
    input [20:0]speed_set_m2;
    input [20:0]speed_set_m3;
    output n20537;
    output n4204;
    output n10;
    output n10_adj_1;
    input VCC_net;
    output n32;
    output n10_adj_2;
    output n10_adj_3;
    output n10_adj_4;
    output n21;
    output n21_adj_5;
    output n21_adj_6;
    output n21_adj_7;
    output n19454;
    output n21_adj_8;
    output n30;
    input \subOut_24__N_1135[1] ;
    input \subOut_24__N_1135[2] ;
    input \subOut_24__N_1135[3] ;
    input \subOut_24__N_1135[4] ;
    input \subOut_24__N_1135[5] ;
    input \subOut_24__N_1135[6] ;
    input \subOut_24__N_1135[7] ;
    input \subOut_24__N_1135[8] ;
    input \subOut_24__N_1135[9] ;
    input \subOut_24__N_1135[10] ;
    input \subOut_24__N_1135[11] ;
    input \subOut_24__N_1135[12] ;
    input \subOut_24__N_1135[13] ;
    input \subOut_24__N_1135[14] ;
    input \subOut_24__N_1135[15] ;
    input \subOut_24__N_1135[16] ;
    input \subOut_24__N_1135[17] ;
    input \subOut_24__N_1135[18] ;
    input \subOut_24__N_1135[19] ;
    input \subOut_24__N_1135[20] ;
    input \subOut_24__N_1135[21] ;
    input \subOut_24__N_1135[24] ;
    input \speed_m1[3] ;
    input [20:0]speed_set_m1;
    input [20:0]speed_set_m4;
    input \speed_m1[7] ;
    input \speed_m1[8] ;
    input \speed_m1[9] ;
    input \speed_m1[12] ;
    input \speed_m1[19] ;
    input \speed_m2[19] ;
    output n5;
    input \speed_m1[1] ;
    input \speed_m2[1] ;
    input \speed_m1[2] ;
    input \speed_m2[2] ;
    input \speed_m1[4] ;
    input \speed_m2[4] ;
    input \speed_m1[5] ;
    input \speed_m2[5] ;
    input \speed_m1[6] ;
    input \speed_m2[6] ;
    input \speed_m1[10] ;
    input \speed_m2[10] ;
    input \speed_m1[11] ;
    input \speed_m2[11] ;
    input \speed_m1[13] ;
    input \speed_m2[13] ;
    input \speed_m1[14] ;
    input \speed_m2[14] ;
    input \speed_m1[15] ;
    input \speed_m2[15] ;
    input \speed_m1[16] ;
    input \speed_m2[16] ;
    input \speed_m1[17] ;
    input \speed_m2[17] ;
    input \speed_m1[18] ;
    input \speed_m2[18] ;
    input \speed_m1[0] ;
    input \speed_m2[0] ;
    output [9:0]PWMdut_m4;
    output [9:0]PWMdut_m3;
    input \speed_m3[3] ;
    input \speed_m2[3] ;
    output n20525;
    input \speed_m3[7] ;
    input \speed_m2[7] ;
    input \speed_m3[8] ;
    input \speed_m2[8] ;
    input \speed_m3[9] ;
    input \speed_m2[9] ;
    input \speed_m3[12] ;
    input \speed_m2[12] ;
    input \speed_m4[1] ;
    input \speed_m3[1] ;
    output n21857;
    input \speed_m4[2] ;
    input \speed_m3[2] ;
    input \speed_m4[4] ;
    input \speed_m3[4] ;
    input \speed_m4[5] ;
    input \speed_m3[5] ;
    input \speed_m4[6] ;
    input \speed_m3[6] ;
    input \speed_m4[10] ;
    input \speed_m3[10] ;
    input \speed_m4[11] ;
    input \speed_m3[11] ;
    input \speed_m4[13] ;
    input \speed_m3[13] ;
    input \speed_m4[14] ;
    input \speed_m3[14] ;
    input \speed_m4[15] ;
    input \speed_m3[15] ;
    input \speed_m4[16] ;
    input \speed_m3[16] ;
    input \speed_m4[17] ;
    input \speed_m3[17] ;
    input \speed_m4[18] ;
    input \speed_m3[18] ;
    input \speed_m4[0] ;
    input \speed_m3[0] ;
    output [9:0]PWMdut_m2;
    output n9;
    output [9:0]PWMdut_m1;
    output n20586;
    input n22383;
    output n4208;
    input n7;
    output n4210;
    output n4209;
    output n4212;
    output n4211;
    output n4214;
    output n4213;
    output n4216;
    output n4215;
    output n4218;
    output n4217;
    output n4220;
    output n4219;
    output n4222;
    output n4221;
    output n4224;
    output n4223;
    output n4226;
    output n4225;
    output n4228;
    output n4227;
    output n4229;
    output n4183;
    output n4182;
    input n13;
    output n4185;
    output n4184;
    input n13_adj_9;
    input n13_adj_10;
    output n4187;
    output n4186;
    input n13_adj_11;
    input n13_adj_12;
    output n4189;
    output n4188;
    input n14;
    output n4191;
    output n4190;
    output n4193;
    output n4192;
    output n4195;
    output n4194;
    output n4197;
    output n4196;
    output n4199;
    output n4198;
    
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(30[4:14])
    wire [4:0]ss;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(96[9:11])
    
    wire n15;
    wire [28:0]backOut0;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(77[9:17])
    
    wire clk_N_683_enable_72;
    wire [28:0]backOut3_28__N_1503;
    wire [28:0]backOut1;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(78[9:17])
    
    wire clk_N_683_enable_40;
    wire [28:0]multOut;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(88[9:16])
    wire [53:0]multOut_28__N_1178;
    
    wire n18755;
    wire [21:0]n2245;
    wire [24:0]subIn2;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(83[9:15])
    
    wire n18756, n18667;
    wire [15:0]n1145;
    wire [9:0]n2153;
    
    wire n18668;
    wire [28:0]intgOut0;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(67[9:17])
    
    wire clk_N_683_enable_100;
    wire [28:0]intgOut0_28__N_735;
    wire [28:0]intgOut1;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(68[9:17])
    
    wire clk_N_683_enable_128;
    wire [28:0]intgOut2;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(69[9:17])
    
    wire clk_N_683_enable_156, clk_N_683_enable_184;
    wire [28:0]Out0;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(72[9:13])
    
    wire clk_N_683_enable_212;
    wire [28:0]Out1;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(73[9:13])
    
    wire clk_N_683_enable_240;
    wire [28:0]Out2;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(74[9:13])
    
    wire clk_N_683_enable_268;
    wire [28:0]Out3;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(75[9:13])
    
    wire clk_N_683_enable_296, clk_N_683_enable_324, clk_N_683_enable_352;
    wire [28:0]addOut;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(92[9:15])
    
    wire n18910;
    wire [24:0]subOut;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(84[9:15])
    wire [28:0]backOut2_28__N_1474;
    wire [28:0]backOut1_28__N_1445;
    
    wire n18909, n3636, n30_c;
    wire [15:0]n1166;
    wire [9:0]n2165;
    wire [9:0]n1302;
    
    wire n14_c, n20197, n18754;
    wire [28:0]Out0_28__N_853;
    
    wire n21897, n22375, clk_N_683_enable_392, subIn1_24__N_1300, dirout_m3_N_1578, 
        subIn1_24__N_1113, dirout_m4_N_1581, n21867, n21868, n21824, 
        n21838;
    wire [23:0]multIn2;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(87[9:16])
    
    wire n4148, n21869, n21894, n21839, n21836, n21834, n22388, 
        n21929, n21928, n21848, n6, n21932, n21888, n21931, n18690, 
        n18691;
    wire [19:0]n3691;
    wire [15:0]n1187;
    
    wire n30_adj_1818, n19129, n13098;
    wire [9:0]n2177;
    wire [9:0]n1346;
    
    wire n21866, n49, n21818, n920;
    wire [28:0]intgOut1_28__N_766;
    
    wire n21821;
    wire [15:0]n1208;
    
    wire n30_adj_1819, n13107, n21849, n21850, n21826, n21862, n56, 
        n16074;
    wire [9:0]n2189;
    wire [9:0]n1390;
    
    wire n57, n42, n5086, n21933, n21858, n18669, n18670, n18666, 
        n16318, n2437, n5138, n18671, n5088, n5084, n5082, n5080, 
        n5078, n5076, n5074, n5072, n5070, n21883, n21892;
    wire [28:0]n588;
    
    wire n5068, mult_29s_25s_0_pp_1_2, mult_29s_25s_0_pp_2_4, mult_29s_25s_0_pp_3_6, 
        mult_29s_25s_0_pp_4_8, mult_29s_25s_0_pp_5_10, mult_29s_25s_0_pp_6_12, 
        mult_29s_25s_0_pp_7_14, mult_29s_25s_0_pp_8_16, mult_29s_25s_0_pp_9_18, 
        mult_29s_25s_0_pp_10_20, mult_29s_25s_0_pp_11_22, mult_29s_25s_0_pp_12_24, 
        mult_29s_25s_0_pp_12_25, mult_29s_25s_0_pp_12_26, mult_29s_25s_0_pp_12_27, 
        mult_29s_25s_0_pp_12_28, mult_29s_25s_0_cin_lr_2, mult_29s_25s_0_cin_lr_4, 
        mult_29s_25s_0_cin_lr_6, mult_29s_25s_0_cin_lr_8, mult_29s_25s_0_cin_lr_10, 
        mult_29s_25s_0_cin_lr_12, mult_29s_25s_0_cin_lr_14, mult_29s_25s_0_cin_lr_16, 
        mult_29s_25s_0_cin_lr_18, mult_29s_25s_0_cin_lr_20, mult_29s_25s_0_cin_lr_22, 
        co_mult_29s_25s_0_0_1, mult_29s_25s_0_pp_0_2, co_mult_29s_25s_0_0_2, 
        s_mult_29s_25s_0_0_4, mult_29s_25s_0_pp_0_4, mult_29s_25s_0_pp_0_3, 
        mult_29s_25s_0_pp_1_4, mult_29s_25s_0_pp_1_3, co_mult_29s_25s_0_0_3, 
        s_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_6, mult_29s_25s_0_pp_0_6, 
        mult_29s_25s_0_pp_0_5, mult_29s_25s_0_pp_1_6, mult_29s_25s_0_pp_1_5, 
        co_mult_29s_25s_0_0_4, s_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_8, 
        mult_29s_25s_0_pp_0_8, mult_29s_25s_0_pp_0_7, mult_29s_25s_0_pp_1_8, 
        mult_29s_25s_0_pp_1_7, co_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_10, mult_29s_25s_0_pp_0_10, mult_29s_25s_0_pp_0_9, 
        mult_29s_25s_0_pp_1_10, mult_29s_25s_0_pp_1_9, co_mult_29s_25s_0_0_6, 
        s_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_12, mult_29s_25s_0_pp_0_12, 
        mult_29s_25s_0_pp_0_11, mult_29s_25s_0_pp_1_12, mult_29s_25s_0_pp_1_11, 
        co_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_14, 
        mult_29s_25s_0_pp_0_14, mult_29s_25s_0_pp_0_13, mult_29s_25s_0_pp_1_14, 
        mult_29s_25s_0_pp_1_13, co_mult_29s_25s_0_0_8, s_mult_29s_25s_0_0_15, 
        s_mult_29s_25s_0_0_16, mult_29s_25s_0_pp_0_16, mult_29s_25s_0_pp_0_15, 
        mult_29s_25s_0_pp_1_16, mult_29s_25s_0_pp_1_15, co_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_17, s_mult_29s_25s_0_0_18, mult_29s_25s_0_pp_0_18, 
        mult_29s_25s_0_pp_0_17, mult_29s_25s_0_pp_1_18, mult_29s_25s_0_pp_1_17, 
        co_mult_29s_25s_0_0_10, s_mult_29s_25s_0_0_19, s_mult_29s_25s_0_0_20, 
        mult_29s_25s_0_pp_0_20, mult_29s_25s_0_pp_0_19, mult_29s_25s_0_pp_1_20, 
        mult_29s_25s_0_pp_1_19, co_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_21, 
        s_mult_29s_25s_0_0_22, mult_29s_25s_0_pp_0_22, mult_29s_25s_0_pp_0_21, 
        mult_29s_25s_0_pp_1_22, mult_29s_25s_0_pp_1_21, co_mult_29s_25s_0_0_12, 
        s_mult_29s_25s_0_0_23, s_mult_29s_25s_0_0_24, mult_29s_25s_0_pp_0_24, 
        mult_29s_25s_0_pp_0_23, mult_29s_25s_0_pp_1_24, mult_29s_25s_0_pp_1_23, 
        co_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_25, s_mult_29s_25s_0_0_26, 
        mult_29s_25s_0_pp_0_26, mult_29s_25s_0_pp_0_25, mult_29s_25s_0_pp_1_26, 
        mult_29s_25s_0_pp_1_25, s_mult_29s_25s_0_0_27, s_mult_29s_25s_0_0_28, 
        mult_29s_25s_0_pp_0_28, mult_29s_25s_0_pp_0_27, mult_29s_25s_0_pp_1_28, 
        mult_29s_25s_0_pp_1_27, co_mult_29s_25s_0_1_1, s_mult_29s_25s_0_1_6, 
        mult_29s_25s_0_pp_2_6, co_mult_29s_25s_0_1_2, s_mult_29s_25s_0_1_7, 
        s_mult_29s_25s_0_1_8, mult_29s_25s_0_pp_2_8, mult_29s_25s_0_pp_2_7, 
        mult_29s_25s_0_pp_3_8, mult_29s_25s_0_pp_3_7, co_mult_29s_25s_0_1_3, 
        s_mult_29s_25s_0_1_9, s_mult_29s_25s_0_1_10, mult_29s_25s_0_pp_2_10, 
        mult_29s_25s_0_pp_2_9, mult_29s_25s_0_pp_3_10, mult_29s_25s_0_pp_3_9, 
        co_mult_29s_25s_0_1_4, s_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_12, 
        mult_29s_25s_0_pp_2_12, mult_29s_25s_0_pp_2_11, mult_29s_25s_0_pp_3_12, 
        mult_29s_25s_0_pp_3_11, co_mult_29s_25s_0_1_5, s_mult_29s_25s_0_1_13, 
        s_mult_29s_25s_0_1_14, mult_29s_25s_0_pp_2_14, mult_29s_25s_0_pp_2_13, 
        mult_29s_25s_0_pp_3_14, mult_29s_25s_0_pp_3_13, co_mult_29s_25s_0_1_6, 
        s_mult_29s_25s_0_1_15, s_mult_29s_25s_0_1_16, mult_29s_25s_0_pp_2_16, 
        mult_29s_25s_0_pp_2_15, mult_29s_25s_0_pp_3_16, mult_29s_25s_0_pp_3_15, 
        co_mult_29s_25s_0_1_7, s_mult_29s_25s_0_1_17, s_mult_29s_25s_0_1_18, 
        mult_29s_25s_0_pp_2_18, mult_29s_25s_0_pp_2_17, mult_29s_25s_0_pp_3_18, 
        mult_29s_25s_0_pp_3_17, co_mult_29s_25s_0_1_8, s_mult_29s_25s_0_1_19, 
        s_mult_29s_25s_0_1_20, mult_29s_25s_0_pp_2_20, mult_29s_25s_0_pp_2_19, 
        mult_29s_25s_0_pp_3_20, mult_29s_25s_0_pp_3_19, co_mult_29s_25s_0_1_9, 
        s_mult_29s_25s_0_1_21, s_mult_29s_25s_0_1_22, mult_29s_25s_0_pp_2_22, 
        mult_29s_25s_0_pp_2_21, mult_29s_25s_0_pp_3_22, mult_29s_25s_0_pp_3_21, 
        co_mult_29s_25s_0_1_10, s_mult_29s_25s_0_1_23, s_mult_29s_25s_0_1_24, 
        mult_29s_25s_0_pp_2_24, mult_29s_25s_0_pp_2_23, mult_29s_25s_0_pp_3_24, 
        mult_29s_25s_0_pp_3_23, co_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_25, 
        s_mult_29s_25s_0_1_26, mult_29s_25s_0_pp_2_26, mult_29s_25s_0_pp_2_25, 
        mult_29s_25s_0_pp_3_26, mult_29s_25s_0_pp_3_25, s_mult_29s_25s_0_1_27, 
        s_mult_29s_25s_0_1_28, mult_29s_25s_0_pp_2_28, mult_29s_25s_0_pp_2_27, 
        mult_29s_25s_0_pp_3_28, mult_29s_25s_0_pp_3_27, co_mult_29s_25s_0_2_1, 
        s_mult_29s_25s_0_2_10, mult_29s_25s_0_pp_4_10, co_mult_29s_25s_0_2_2, 
        s_mult_29s_25s_0_2_12, s_mult_29s_25s_0_2_11, mult_29s_25s_0_pp_4_12, 
        mult_29s_25s_0_pp_4_11, mult_29s_25s_0_pp_5_12, mult_29s_25s_0_pp_5_11, 
        co_mult_29s_25s_0_2_3, s_mult_29s_25s_0_2_13, s_mult_29s_25s_0_2_14, 
        mult_29s_25s_0_pp_4_14, mult_29s_25s_0_pp_4_13, mult_29s_25s_0_pp_5_14, 
        mult_29s_25s_0_pp_5_13, co_mult_29s_25s_0_2_4, s_mult_29s_25s_0_2_15, 
        s_mult_29s_25s_0_2_16, mult_29s_25s_0_pp_4_16, mult_29s_25s_0_pp_4_15, 
        mult_29s_25s_0_pp_5_16, mult_29s_25s_0_pp_5_15, co_mult_29s_25s_0_2_5, 
        s_mult_29s_25s_0_2_17, s_mult_29s_25s_0_2_18, mult_29s_25s_0_pp_4_18, 
        mult_29s_25s_0_pp_4_17, mult_29s_25s_0_pp_5_18, mult_29s_25s_0_pp_5_17, 
        co_mult_29s_25s_0_2_6, s_mult_29s_25s_0_2_19, s_mult_29s_25s_0_2_20, 
        mult_29s_25s_0_pp_4_20, mult_29s_25s_0_pp_4_19, mult_29s_25s_0_pp_5_20, 
        mult_29s_25s_0_pp_5_19, co_mult_29s_25s_0_2_7, s_mult_29s_25s_0_2_21, 
        s_mult_29s_25s_0_2_22, mult_29s_25s_0_pp_4_22, mult_29s_25s_0_pp_4_21, 
        mult_29s_25s_0_pp_5_22, mult_29s_25s_0_pp_5_21, co_mult_29s_25s_0_2_8, 
        s_mult_29s_25s_0_2_23, s_mult_29s_25s_0_2_24, mult_29s_25s_0_pp_4_24, 
        mult_29s_25s_0_pp_4_23, mult_29s_25s_0_pp_5_24, mult_29s_25s_0_pp_5_23, 
        co_mult_29s_25s_0_2_9, s_mult_29s_25s_0_2_25, s_mult_29s_25s_0_2_26, 
        mult_29s_25s_0_pp_4_26, mult_29s_25s_0_pp_4_25, mult_29s_25s_0_pp_5_26, 
        mult_29s_25s_0_pp_5_25, s_mult_29s_25s_0_2_27, s_mult_29s_25s_0_2_28, 
        mult_29s_25s_0_pp_4_28, mult_29s_25s_0_pp_4_27, mult_29s_25s_0_pp_5_28, 
        mult_29s_25s_0_pp_5_27, co_mult_29s_25s_0_3_1, s_mult_29s_25s_0_3_14, 
        mult_29s_25s_0_pp_6_14, co_mult_29s_25s_0_3_2, s_mult_29s_25s_0_3_15, 
        s_mult_29s_25s_0_3_16, mult_29s_25s_0_pp_6_16, mult_29s_25s_0_pp_6_15, 
        mult_29s_25s_0_pp_7_16, mult_29s_25s_0_pp_7_15, co_mult_29s_25s_0_3_3, 
        s_mult_29s_25s_0_3_17, s_mult_29s_25s_0_3_18, mult_29s_25s_0_pp_6_18, 
        mult_29s_25s_0_pp_6_17, mult_29s_25s_0_pp_7_18, mult_29s_25s_0_pp_7_17, 
        co_mult_29s_25s_0_3_4, s_mult_29s_25s_0_3_19, s_mult_29s_25s_0_3_20, 
        mult_29s_25s_0_pp_6_20, mult_29s_25s_0_pp_6_19, mult_29s_25s_0_pp_7_20, 
        mult_29s_25s_0_pp_7_19, co_mult_29s_25s_0_3_5, s_mult_29s_25s_0_3_21, 
        s_mult_29s_25s_0_3_22, mult_29s_25s_0_pp_6_22, mult_29s_25s_0_pp_6_21, 
        mult_29s_25s_0_pp_7_22, mult_29s_25s_0_pp_7_21, co_mult_29s_25s_0_3_6, 
        s_mult_29s_25s_0_3_23, s_mult_29s_25s_0_3_24, mult_29s_25s_0_pp_6_24, 
        mult_29s_25s_0_pp_6_23, mult_29s_25s_0_pp_7_24, mult_29s_25s_0_pp_7_23, 
        co_mult_29s_25s_0_3_7, s_mult_29s_25s_0_3_25, s_mult_29s_25s_0_3_26, 
        mult_29s_25s_0_pp_6_26, mult_29s_25s_0_pp_6_25, mult_29s_25s_0_pp_7_26, 
        mult_29s_25s_0_pp_7_25, s_mult_29s_25s_0_3_27, s_mult_29s_25s_0_3_28, 
        mult_29s_25s_0_pp_6_28, mult_29s_25s_0_pp_6_27, mult_29s_25s_0_pp_7_28, 
        mult_29s_25s_0_pp_7_27, co_mult_29s_25s_0_4_1, s_mult_29s_25s_0_4_18, 
        mult_29s_25s_0_pp_8_18, co_mult_29s_25s_0_4_2, s_mult_29s_25s_0_4_20, 
        s_mult_29s_25s_0_4_19, mult_29s_25s_0_pp_8_20, mult_29s_25s_0_pp_8_19, 
        mult_29s_25s_0_pp_9_20, mult_29s_25s_0_pp_9_19, co_mult_29s_25s_0_4_3, 
        s_mult_29s_25s_0_4_21, s_mult_29s_25s_0_4_22, mult_29s_25s_0_pp_8_22, 
        mult_29s_25s_0_pp_8_21, mult_29s_25s_0_pp_9_22, mult_29s_25s_0_pp_9_21, 
        co_mult_29s_25s_0_4_4, s_mult_29s_25s_0_4_23, s_mult_29s_25s_0_4_24, 
        mult_29s_25s_0_pp_8_24, mult_29s_25s_0_pp_8_23, mult_29s_25s_0_pp_9_24, 
        mult_29s_25s_0_pp_9_23, co_mult_29s_25s_0_4_5, s_mult_29s_25s_0_4_25, 
        s_mult_29s_25s_0_4_26, mult_29s_25s_0_pp_8_26, mult_29s_25s_0_pp_8_25, 
        mult_29s_25s_0_pp_9_26, mult_29s_25s_0_pp_9_25, s_mult_29s_25s_0_4_27, 
        s_mult_29s_25s_0_4_28, mult_29s_25s_0_pp_8_28, mult_29s_25s_0_pp_8_27, 
        mult_29s_25s_0_pp_9_28, mult_29s_25s_0_pp_9_27, co_mult_29s_25s_0_5_1, 
        s_mult_29s_25s_0_5_22, mult_29s_25s_0_pp_10_22, co_mult_29s_25s_0_5_2, 
        s_mult_29s_25s_0_5_23, s_mult_29s_25s_0_5_24, mult_29s_25s_0_pp_10_24, 
        mult_29s_25s_0_pp_10_23, mult_29s_25s_0_pp_11_24, mult_29s_25s_0_pp_11_23, 
        co_mult_29s_25s_0_5_3, s_mult_29s_25s_0_5_25, s_mult_29s_25s_0_5_26, 
        mult_29s_25s_0_pp_10_26, mult_29s_25s_0_pp_10_25, mult_29s_25s_0_pp_11_26, 
        mult_29s_25s_0_pp_11_25, s_mult_29s_25s_0_5_27, s_mult_29s_25s_0_5_28, 
        mult_29s_25s_0_pp_10_28, mult_29s_25s_0_pp_10_27, mult_29s_25s_0_pp_11_28, 
        mult_29s_25s_0_pp_11_27, co_mult_29s_25s_0_6_1, s_mult_29s_25s_0_6_24, 
        co_mult_29s_25s_0_6_2, s_mult_29s_25s_0_6_25, s_mult_29s_25s_0_6_26, 
        s_mult_29s_25s_0_6_27, s_mult_29s_25s_0_6_28, co_mult_29s_25s_0_7_1, 
        co_mult_29s_25s_0_7_2, mult_29s_25s_0_pp_2_5, co_mult_29s_25s_0_7_3, 
        s_mult_29s_25s_0_7_8, co_mult_29s_25s_0_7_4, s_mult_29s_25s_0_7_9, 
        s_mult_29s_25s_0_7_10, co_mult_29s_25s_0_7_5, s_mult_29s_25s_0_7_11, 
        s_mult_29s_25s_0_7_12, co_mult_29s_25s_0_7_6, s_mult_29s_25s_0_7_13, 
        s_mult_29s_25s_0_7_14, co_mult_29s_25s_0_7_7, s_mult_29s_25s_0_7_15, 
        s_mult_29s_25s_0_7_16, co_mult_29s_25s_0_7_8, s_mult_29s_25s_0_7_17, 
        s_mult_29s_25s_0_7_18, co_mult_29s_25s_0_7_9, s_mult_29s_25s_0_7_19, 
        s_mult_29s_25s_0_7_20, co_mult_29s_25s_0_7_10, s_mult_29s_25s_0_7_21, 
        s_mult_29s_25s_0_7_22, co_mult_29s_25s_0_7_11, s_mult_29s_25s_0_7_23, 
        s_mult_29s_25s_0_7_24, co_mult_29s_25s_0_7_12, s_mult_29s_25s_0_7_25, 
        s_mult_29s_25s_0_7_26, s_mult_29s_25s_0_7_27, s_mult_29s_25s_0_7_28, 
        n5066, co_mult_29s_25s_0_8_1, s_mult_29s_25s_0_8_12, co_mult_29s_25s_0_8_2, 
        s_mult_29s_25s_0_8_13, s_mult_29s_25s_0_8_14, mult_29s_25s_0_pp_6_13, 
        co_mult_29s_25s_0_8_3, s_mult_29s_25s_0_8_15, s_mult_29s_25s_0_8_16, 
        co_mult_29s_25s_0_8_4, s_mult_29s_25s_0_8_17, s_mult_29s_25s_0_8_18, 
        co_mult_29s_25s_0_8_5, s_mult_29s_25s_0_8_19, s_mult_29s_25s_0_8_20, 
        co_mult_29s_25s_0_8_6, s_mult_29s_25s_0_8_21, s_mult_29s_25s_0_8_22, 
        co_mult_29s_25s_0_8_7, s_mult_29s_25s_0_8_23, s_mult_29s_25s_0_8_24, 
        co_mult_29s_25s_0_8_8, s_mult_29s_25s_0_8_25, s_mult_29s_25s_0_8_26, 
        s_mult_29s_25s_0_8_27, s_mult_29s_25s_0_8_28, n21926, n5064, 
        co_mult_29s_25s_0_9_1, s_mult_29s_25s_0_9_20, co_mult_29s_25s_0_9_2, 
        s_mult_29s_25s_0_9_21, s_mult_29s_25s_0_9_22, mult_29s_25s_0_pp_10_21, 
        co_mult_29s_25s_0_9_3, s_mult_29s_25s_0_9_24, s_mult_29s_25s_0_9_23, 
        co_mult_29s_25s_0_9_4, s_mult_29s_25s_0_9_25, s_mult_29s_25s_0_9_26, 
        s_mult_29s_25s_0_9_27, s_mult_29s_25s_0_9_28, co_mult_29s_25s_0_10_1, 
        co_mult_29s_25s_0_10_2, mult_29s_25s_0_pp_4_9, co_mult_29s_25s_0_10_3, 
        co_mult_29s_25s_0_10_4, co_mult_29s_25s_0_10_5, s_mult_29s_25s_0_10_16, 
        co_mult_29s_25s_0_10_6, s_mult_29s_25s_0_10_17, s_mult_29s_25s_0_10_18, 
        co_mult_29s_25s_0_10_7, s_mult_29s_25s_0_10_19, s_mult_29s_25s_0_10_20, 
        co_mult_29s_25s_0_10_8, s_mult_29s_25s_0_10_21, s_mult_29s_25s_0_10_22, 
        co_mult_29s_25s_0_10_9, s_mult_29s_25s_0_10_23, s_mult_29s_25s_0_10_24, 
        co_mult_29s_25s_0_10_10, s_mult_29s_25s_0_10_25, s_mult_29s_25s_0_10_26, 
        s_mult_29s_25s_0_10_27, s_mult_29s_25s_0_10_28, n5062, n5060, 
        co_mult_29s_25s_0_11_1, s_mult_29s_25s_0_11_24, co_mult_29s_25s_0_11_2, 
        s_mult_29s_25s_0_11_25, s_mult_29s_25s_0_11_26, s_mult_29s_25s_0_11_27, 
        s_mult_29s_25s_0_11_28, n21884, co_t_mult_29s_25s_0_12_1, co_t_mult_29s_25s_0_12_2, 
        mult_29s_25s_0_pp_8_17, co_t_mult_29s_25s_0_12_3, co_t_mult_29s_25s_0_12_4, 
        co_t_mult_29s_25s_0_12_5, co_t_mult_29s_25s_0_12_6, mult_29s_25s_0_cin_lr_0, 
        mco, mco_1, mco_2, mco_3, mco_4, mco_5, mco_6, mco_7, 
        mco_8, mco_9, mco_10, mco_11, mco_12, mco_14, mco_15, 
        mco_16, mco_17, mco_18, mco_19, mco_20, mco_21, mco_22, 
        mco_23, mco_24, mco_25, mco_28, mco_29, mco_30, mco_31, 
        mco_32, mco_33, mco_34, mco_35, mco_36, mco_37, mco_38, 
        mco_42, mco_43, mco_44, mco_45, mco_46, mco_47, mco_48, 
        mco_49, mco_50, mco_51, mco_56, mco_57, mco_58, mco_59, 
        mco_60, mco_61, mco_62, mco_63, mco_64, mco_70, mco_71, 
        mco_72, mco_73, mco_74, mco_75, mco_76, mco_77, mco_84, 
        mco_85, mco_86, mco_87, mco_88, mco_89, mco_90, mco_98, 
        mco_99, mco_100, mco_101, mco_102, mco_103, mco_112, mco_113, 
        mco_114, mco_115, mco_116, mco_126, mco_127, mco_128, mco_129, 
        mco_140, mco_141, mco_142, mco_154, mco_155, n5058, n14_adj_1824, 
        n10_adj_1825, n19130, n20184, n6_adj_1826, n19131;
    wire [28:0]n121;
    
    wire n5056, n5054, n21820, n21925;
    wire [28:0]n648;
    wire [28:0]n678;
    
    wire n18908, n19086, n19087, n21817, n5052, n5050, n23, n23_adj_1827, 
        n23_adj_1829, n23_adj_1831, n18907, n21815, n7_c;
    wire [28:0]intgOut2_28__N_795;
    wire [28:0]intgOut3_c;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(70[9:17])
    wire [28:0]backOut2_c;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(79[9:17])
    wire [28:0]backOut3_c;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(80[9:17])
    
    wire n23_adj_1833, n28, n21870, n5046, n16214, n21816, n21877;
    wire [20:0]subIn2_24__N_1301;
    wire [20:0]subIn2_24__N_1114;
    
    wire n35, n5100, n5122, n5128, n5124, n9_c, n7_adj_1836, n18906, 
        n10_adj_1837, n8, n4, n5118, n5098, n5108, n5114, n18905, 
        n18904, n9_adj_1838, n7_adj_1839, n10_adj_1840, n8_adj_1841, 
        n4_adj_1842, n5110, n5106, n18689, n5104, n5102, n18903, 
        n5048, n5092, n5126, n13082, n18688, n5116, n5096, n22376, 
        n5094, n5120, n5130, n21885, n20247, n21903, n5112, n20202, 
        n20199, n9_adj_1843, n7_adj_1844, n10_adj_1845, n8_adj_1846, 
        n4_adj_1847;
    wire [21:0]n2485;
    
    wire n18902, n18901, n18900, n16286;
    wire [28:0]n558;
    
    wire n18899, n13089, n13080;
    wire [9:0]n1258;
    
    wire n5707, n18687, n5689, n5691, n5693, n5695, n5697, n18898, 
        n18686, n21819, n5699, n5701, n9_adj_1849, n7_adj_1850, 
        n30_adj_1851, n10_adj_1852, n18897, n8_adj_1853, n4_adj_1854, 
        n5703, n18896, n14_adj_1855, n10_adj_1856, n19124, n6_adj_1857, 
        n19125, n21922, n21898, n21893, n5705, n22379, n5709, 
        n5711, n18685, n21923, n21886, n5713, n5715, n18684, n18683, 
        n5717, n18682, n5719, n5721, n5723, n5725, n18681, n5178, 
        n18878, n18877, n5729, n18680, n5176, n18876, n18679, 
        n5172, n5174, n18875, n5254, n18874, n20055, n18991, n18990, 
        n21924, n18678, n5168, n5170, n18989, n18988, n18987, 
        n18986, n18985, n18873, n18872, n18984, n18780, n18983, 
        n18871, n18982, n18981, n18980, n18677, n5164, n5166, 
        n18979, n18779, n18978, n18977, n18976, n18870, n5162, 
        n5160, n18975, n5158, n5156, n18974, n18869, n18973, n18972, 
        n5154, n5152, n5150, n5148, n5146, n5144, n5142, n5140, 
        n5690, n5692, n5694, n5696, n5698, n5700, n18868, n5702, 
        n5704, n5706, n5708, n18867, n5710, n18866, n5712, n5714, 
        n5716, n5718, n18865, n5720, n5722, n5724, n18864, n18863, 
        n5726, n5730, n5255, n18862, n18861;
    wire [28:0]n618;
    wire [28:0]addIn2_28__N_1337;
    wire [28:0]addIn2_28__N_1207;
    
    wire n18860, n18859, n14_adj_1858, n10_adj_1859, n20582, n18858, 
        n6_adj_1860, n18857, n18778, n18777, n18856, n18855, n18854, 
        n18853, n18852, n18851, n18776, n18850, n18849, n18676, 
        n18848, n21895, n18775, n18713, n18774, n18712, n18675, 
        n18773, n18711, n18772, n18710, n18674, n18673, n14_adj_1862, 
        n10_adj_1863, n19127, n6_adj_1864, n19128, n18771, n18709, 
        n18708, n18707, n18706, n18834, n18770, n18672, n18833, 
        n18705, n18832, n18920, n18919, n18831, n18769, n18704, 
        n18830, n18918, n18703, n18829, n18828, n18768, n18702, 
        n18827, n18917, n18767, n18701, n18826, n18916, n18700, 
        n18766, n18825, n18699, n18824, n18915, n18764, n18698, 
        n18823, n18914, n18763, n18822, n18762, n18697, n18821, 
        n18913, n18761, n18696, n18912, n18695, n18760, n18759, 
        n18694, n18911, n18758, n18693, n18692, n18757;
    
    LUT4 i8798_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[2]), .C(ss[3]), .D(ss[1]), 
         .Z(n15)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i8798_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3AX backOut0_i0_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i0.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i0.GSR = "DISABLED";
    FD1S3AX multOut_i0 (.D(multOut_28__N_1178[0]), .CK(clk_N_683), .Q(multOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i0.GSR = "ENABLED";
    CCU2D sub_17_rep_2_add_2_5 (.A0(n2245[3]), .B0(subIn2[3]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[4]), .B1(subIn2[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18755), .COUT(n18756), .S0(n4201), .S1(n4200));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_5.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_5.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_5.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_5.INJECT1_1 = "NO";
    CCU2D add_1174_5 (.A0(n1145[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18667), 
          .COUT(n18668), .S0(n2153[3]), .S1(n2153[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(327[20:29])
    defparam add_1174_5.INIT0 = 16'hf555;
    defparam add_1174_5.INIT1 = 16'hf555;
    defparam add_1174_5.INJECT1_0 = "NO";
    defparam add_1174_5.INJECT1_1 = "NO";
    FD1P3AX intgOut0_i0 (.D(intgOut0_28__N_735[0]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i0.GSR = "ENABLED";
    FD1P3AX intgOut1_i0 (.D(intgOut0_28__N_735[0]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i0.GSR = "ENABLED";
    FD1P3AX intgOut2_i0 (.D(intgOut0_28__N_735[0]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i0.GSR = "ENABLED";
    FD1P3AX intgOut3_i0 (.D(intgOut0_28__N_735[0]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i0.GSR = "ENABLED";
    FD1P3AX Out0_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i0.GSR = "ENABLED";
    FD1P3AX Out1_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i0.GSR = "ENABLED";
    FD1P3AX Out2_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i0.GSR = "ENABLED";
    FD1P3AX Out3_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i0.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i0.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i0 (.D(backOut3_28__N_1503[0]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i0.GSR = "DISABLED";
    CCU2D add_16119_2 (.A0(addOut[7]), .B0(addOut[6]), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18910));
    defparam add_16119_2.INIT0 = 16'h1000;
    defparam add_16119_2.INIT1 = 16'h5555;
    defparam add_16119_2.INJECT1_0 = "NO";
    defparam add_16119_2.INJECT1_1 = "NO";
    FD1S3AX subOut_i0 (.D(\subOut_24__N_1135[0] ), .CK(clk_N_683), .Q(subOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i0.GSR = "ENABLED";
    FD1P3AX backOut1_i0_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i23.GSR = "DISABLED";
    CCU2D add_16120_29 (.A0(addOut[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18909), 
          .S1(n3636));
    defparam add_16120_29.INIT0 = 16'h5aaa;
    defparam add_16120_29.INIT1 = 16'h0000;
    defparam add_16120_29.INJECT1_0 = "NO";
    defparam add_16120_29.INJECT1_1 = "NO";
    FD1P3AX backOut1_i0_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i22.GSR = "DISABLED";
    LUT4 mux_205_i9_3_lut_4_lut_3_lut (.A(n30_c), .B(n1166[15]), .C(n2165[8]), 
         .Z(n1302[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(334[25:42])
    defparam mux_205_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FD1P3AX backOut1_i0_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i13.GSR = "DISABLED";
    FD1S3IX ss_i2 (.D(n14_c), .CK(clk_N_683), .CD(ss[4]), .Q(ss[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam ss_i2.GSR = "ENABLED";
    FD1S3IX ss_i3 (.D(n15), .CK(clk_N_683), .CD(ss[4]), .Q(ss[3]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam ss_i3.GSR = "ENABLED";
    FD1S3AY ss_i4 (.D(n20197), .CK(clk_N_683), .Q(ss[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam ss_i4.GSR = "ENABLED";
    FD1P3AX backOut1_i0_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i11.GSR = "DISABLED";
    CCU2D sub_17_rep_2_add_2_3 (.A0(n2245[1]), .B0(subIn2[1]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[2]), .B1(subIn2[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18754), .COUT(n18755), .S0(n4203), .S1(n4202));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_3.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_3.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_3.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_3.INJECT1_1 = "NO";
    FD1P3AX backOut1_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_40), 
            .CK(clk_N_683), .Q(backOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i1.GSR = "DISABLED";
    FD1S3IX ss_i0 (.D(n21897), .CK(clk_N_683), .CD(ss[4]), .Q(ss[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam ss_i0.GSR = "ENABLED";
    FD1S3IX ss_i1 (.D(n22375), .CK(clk_N_683), .CD(ss[4]), .Q(ss[1]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam ss_i1.GSR = "ENABLED";
    FD1P3AX dirout_m2_308 (.D(subIn1_24__N_1300), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m2));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dirout_m2_308.GSR = "DISABLED";
    FD1P3AX dirout_m3_309 (.D(dirout_m3_N_1578), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m3));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dirout_m3_309.GSR = "DISABLED";
    FD1P3AX dirout_m1_307 (.D(subIn1_24__N_1113), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m1));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dirout_m1_307.GSR = "DISABLED";
    FD1P3AX dirout_m4_310 (.D(dirout_m4_N_1581), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m4));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dirout_m4_310.GSR = "DISABLED";
    LUT4 i13973_3_lut_rep_404_3_lut_4_lut_4_lut_4_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21867), .D(n21868), .Z(n21824)) /* synthesis lut_function=(A (B+(C (D)))+!A ((C)+!B)) */ ;
    defparam i13973_3_lut_rep_404_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hf9d9;
    LUT4 i13240_3_lut_4_lut (.A(n21851), .B(n21838), .C(multIn2[6]), .D(n4148), 
         .Z(multIn2[3])) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i13240_3_lut_4_lut.init = 16'hff07;
    LUT4 ss_2__bdd_3_lut_rep_419_4_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21869), 
         .D(n21894), .Z(n21839)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(170[9:16])
    defparam ss_2__bdd_3_lut_rep_419_4_lut_4_lut.init = 16'hf7e6;
    LUT4 i1_3_lut_rep_416_4_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21868), 
         .D(n21869), .Z(n21836)) /* synthesis lut_function=(A+(B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(172[20:27])
    defparam i1_3_lut_rep_416_4_lut_4_lut.init = 16'hfbea;
    LUT4 i2_3_lut_rep_414_4_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21868), 
         .D(n21869), .Z(n21834)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((D)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam i2_3_lut_rep_414_4_lut_4_lut.init = 16'hf791;
    LUT4 i13239_3_lut_4_lut (.A(n21851), .B(n21838), .C(multIn2[6]), .D(n4148), 
         .Z(multIn2[5])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;
    defparam i13239_3_lut_4_lut.init = 16'h00f7;
    LUT4 i1_4_lut_then_4_lut (.A(n22388), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21929)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_else_4_lut (.A(n22388), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21928)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0100;
    LUT4 i1839_2_lut_rep_505 (.A(ss[0]), .B(ss[1]), .Z(n22375)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1839_2_lut_rep_505.init = 16'h6666;
    LUT4 i18047_3_lut_3_lut_4_lut_4_lut_then_4_lut (.A(ss[3]), .B(n22388), 
         .C(n21848), .D(n6), .Z(n21932)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam i18047_3_lut_3_lut_4_lut_4_lut_then_4_lut.init = 16'hf0d0;
    LUT4 i18047_3_lut_3_lut_4_lut_4_lut_else_4_lut (.A(ss[3]), .B(n22388), 
         .C(n21848), .D(n21888), .Z(n21931)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam i18047_3_lut_3_lut_4_lut_4_lut_else_4_lut.init = 16'hf0d0;
    LUT4 mux_205_i10_3_lut_4_lut_3_lut (.A(n30_c), .B(n1166[15]), .C(n2165[9]), 
         .Z(n1302[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(334[25:42])
    defparam mux_205_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    CCU2D add_183_3 (.A0(Out1[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18690), 
          .COUT(n18691), .S0(n1166[1]), .S1(n1166[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_3.INIT0 = 16'h5aaa;
    defparam add_183_3.INIT1 = 16'h5aaa;
    defparam add_183_3.INJECT1_0 = "NO";
    defparam add_183_3.INJECT1_1 = "NO";
    LUT4 mux_205_i8_3_lut_4_lut_3_lut (.A(n30_c), .B(n1166[15]), .C(n2165[7]), 
         .Z(n1302[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(334[25:42])
    defparam mux_205_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_205_i6_3_lut_4_lut_3_lut (.A(n30_c), .B(n1166[15]), .C(n2165[5]), 
         .Z(n1302[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(334[25:42])
    defparam mux_205_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_1799_i4_3_lut_4_lut_4_lut (.A(n21835), .B(\speed_m4[3] ), .C(n4133), 
         .D(n21838), .Z(n3691[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam mux_1799_i4_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 i10668_3_lut_4_lut (.A(n1187[15]), .B(n30_adj_1818), .C(n19129), 
         .D(clk_N_683_enable_392), .Z(n13098)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(342[7:42])
    defparam i10668_3_lut_4_lut.init = 16'hf700;
    LUT4 mux_1799_i8_3_lut_4_lut_4_lut (.A(n21835), .B(\speed_m4[7] ), .C(n4133), 
         .D(n21838), .Z(n3691[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam mux_1799_i8_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_1799_i9_3_lut_4_lut_4_lut (.A(n21835), .B(\speed_m4[8] ), .C(n4133), 
         .D(n21838), .Z(n3691[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam mux_1799_i9_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_1799_i10_3_lut_4_lut_4_lut (.A(n21835), .B(\speed_m4[9] ), 
         .C(n4133), .D(n21838), .Z(n3691[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam mux_1799_i10_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_1799_i13_3_lut_4_lut_4_lut (.A(n21835), .B(\speed_m4[12] ), 
         .C(n4133), .D(n21838), .Z(n3691[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam mux_1799_i13_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_212_i4_3_lut_4_lut_3_lut (.A(n30_adj_1818), .B(n1187[15]), 
         .C(n2177[3]), .Z(n1346[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(342[25:42])
    defparam mux_212_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i52_2_lut_rep_398_4_lut (.A(n21848), .B(n21869), .C(n21866), 
         .D(n49), .Z(n21818)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(D))) */ ;
    defparam i52_2_lut_rep_398_4_lut.init = 16'h5700;
    LUT4 mux_212_i10_3_lut_4_lut_3_lut (.A(n30_adj_1818), .B(n1187[15]), 
         .C(n2177[9]), .Z(n1346[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(342[25:42])
    defparam mux_212_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FD1S3AY ss_i4_rep_516 (.D(n20197), .CK(clk_N_683), .Q(n22388));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam ss_i4_rep_516.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n920), .B(n3636), .C(addOut[1]), .D(n22388), 
         .Z(intgOut1_28__N_766[1])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_212_i7_3_lut_4_lut_3_lut (.A(n30_adj_1818), .B(n1187[15]), 
         .C(n2177[6]), .Z(n1346[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(342[25:42])
    defparam mux_212_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_212_i9_3_lut_4_lut_3_lut (.A(n30_adj_1818), .B(n1187[15]), 
         .C(n2177[8]), .Z(n1346[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(342[25:42])
    defparam mux_212_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i13815_2_lut_rep_401_4_lut (.A(n21848), .B(n21869), .C(n21866), 
         .D(n49), .Z(n21821)) /* synthesis lut_function=(A (B+(C+(D)))+!A (D)) */ ;
    defparam i13815_2_lut_rep_401_4_lut.init = 16'hffa8;
    LUT4 i13570_4_lut_4_lut (.A(n920), .B(n3636), .C(addOut[14]), .D(n22388), 
         .Z(intgOut1_28__N_766[14])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13570_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_212_i8_3_lut_4_lut_3_lut (.A(n30_adj_1818), .B(n1187[15]), 
         .C(n2177[7]), .Z(n1346[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(342[25:42])
    defparam mux_212_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_212_i6_3_lut_4_lut_3_lut (.A(n30_adj_1818), .B(n1187[15]), 
         .C(n2177[5]), .Z(n1346[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(342[25:42])
    defparam mux_212_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i10670_3_lut_4_lut (.A(n1208[15]), .B(n30_adj_1819), .C(n19129), 
         .D(clk_N_683_enable_392), .Z(n13107)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(350[7:42])
    defparam i10670_3_lut_4_lut.init = 16'hf700;
    LUT4 i1_2_lut_rep_406_4_lut (.A(n21849), .B(n6), .C(n21869), .D(n21850), 
         .Z(n21826)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_406_4_lut.init = 16'ha800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_36 (.A(n920), .B(n3636), .C(addOut[2]), 
         .D(n22388), .Z(intgOut0_28__N_735[2])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_36.init = 16'h0010;
    LUT4 i13817_2_lut_4_lut (.A(n21862), .B(n6), .C(n21894), .D(n56), 
         .Z(n16074)) /* synthesis lut_function=(A (B+(C+(D)))+!A (D)) */ ;
    defparam i13817_2_lut_4_lut.init = 16'hffa8;
    LUT4 mux_219_i4_3_lut_4_lut_3_lut (.A(n30_adj_1819), .B(n1208[15]), 
         .C(n2189[3]), .Z(n1390[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(350[25:42])
    defparam mux_219_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i59_2_lut_4_lut (.A(n21862), .B(n6), .C(n21894), .D(n56), .Z(n57)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(D))) */ ;
    defparam i59_2_lut_4_lut.init = 16'h5700;
    LUT4 mux_219_i10_3_lut_4_lut_3_lut (.A(n30_adj_1819), .B(n1208[15]), 
         .C(n2189[9]), .Z(n1390[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(350[25:42])
    defparam mux_219_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_219_i7_3_lut_4_lut_3_lut (.A(n30_adj_1819), .B(n1208[15]), 
         .C(n2189[6]), .Z(n1390[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(350[25:42])
    defparam mux_219_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i13571_4_lut_4_lut (.A(n920), .B(n3636), .C(addOut[16]), .D(n22388), 
         .Z(intgOut1_28__N_766[16])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13571_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_219_i9_3_lut_4_lut_3_lut (.A(n30_adj_1819), .B(n1208[15]), 
         .C(n2189[8]), .Z(n1390[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(350[25:42])
    defparam mux_219_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_219_i8_3_lut_4_lut_3_lut (.A(n30_adj_1819), .B(n1208[15]), 
         .C(n2189[7]), .Z(n1390[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(350[25:42])
    defparam mux_219_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_219_i6_3_lut_4_lut_3_lut (.A(n30_adj_1819), .B(n1208[15]), 
         .C(n2189[5]), .Z(n1390[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(350[25:42])
    defparam mux_219_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_1190_i20_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[19]), 
         .D(speed_set_m3[19]), .Z(n5086)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_3_lut_4_lut_adj_37 (.A(n920), .B(n3636), .C(addOut[3]), 
         .D(n22388), .Z(intgOut1_28__N_766[3])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_37.init = 16'h0010;
    LUT4 i18348_4_lut_4_lut (.A(n21850), .B(n21933), .C(n21862), .D(n21858), 
         .Z(n20537)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 185[26])
    defparam i18348_4_lut_4_lut.init = 16'hdfff;
    CCU2D add_1174_9 (.A0(n1145[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18669), 
          .COUT(n18670), .S0(n2153[7]), .S1(n2153[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(327[20:29])
    defparam add_1174_9.INIT0 = 16'hf555;
    defparam add_1174_9.INIT1 = 16'hf555;
    defparam add_1174_9.INJECT1_0 = "NO";
    defparam add_1174_9.INJECT1_1 = "NO";
    CCU2D add_1174_3 (.A0(n1145[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18666), 
          .COUT(n18667), .S0(n2153[1]), .S1(n2153[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(327[20:29])
    defparam add_1174_3.INIT0 = 16'hf555;
    defparam add_1174_3.INIT1 = 16'hf555;
    defparam add_1174_3.INJECT1_0 = "NO";
    defparam add_1174_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_38 (.A(n21826), .B(n42), .C(n16318), 
         .D(n21818), .Z(n2437)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam i1_2_lut_3_lut_4_lut_adj_38.init = 16'hf040;
    CCU2D add_1180_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5138), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18671), 
          .S1(n2245[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_1.INIT0 = 16'hF000;
    defparam add_1180_1.INIT1 = 16'h0aaa;
    defparam add_1180_1.INJECT1_0 = "NO";
    defparam add_1180_1.INJECT1_1 = "NO";
    CCU2D add_1174_7 (.A0(n1145[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18668), 
          .COUT(n18669), .S0(n2153[5]), .S1(n2153[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(327[20:29])
    defparam add_1174_7.INIT0 = 16'hf555;
    defparam add_1174_7.INIT1 = 16'hf555;
    defparam add_1174_7.INJECT1_0 = "NO";
    defparam add_1174_7.INJECT1_1 = "NO";
    CCU2D add_1174_11 (.A0(n1145[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18670), 
          .S0(n2153[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(327[20:29])
    defparam add_1174_11.INIT0 = 16'hf555;
    defparam add_1174_11.INIT1 = 16'h0000;
    defparam add_1174_11.INJECT1_0 = "NO";
    defparam add_1174_11.INJECT1_1 = "NO";
    CCU2D add_1174_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18666), 
          .S1(n2153[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(327[20:29])
    defparam add_1174_1.INIT0 = 16'hF000;
    defparam add_1174_1.INIT1 = 16'h0aaa;
    defparam add_1174_1.INJECT1_0 = "NO";
    defparam add_1174_1.INJECT1_1 = "NO";
    LUT4 mux_1190_i21_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[20]), 
         .D(speed_set_m3[20]), .Z(n5088)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i19_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[18]), 
         .D(speed_set_m3[18]), .Z(n5084)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i18_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[17]), 
         .D(speed_set_m3[17]), .Z(n5082)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i17_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[16]), 
         .D(speed_set_m3[16]), .Z(n5080)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i16_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[15]), 
         .D(speed_set_m3[15]), .Z(n5078)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i15_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[14]), 
         .D(speed_set_m3[14]), .Z(n5076)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i14_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[13]), 
         .D(speed_set_m3[13]), .Z(n5074)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i13_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[12]), 
         .D(speed_set_m3[12]), .Z(n5072)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i12_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[11]), 
         .D(speed_set_m3[11]), .Z(n5070)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13563_4_lut_4_lut (.A(n920), .B(n3636), .C(addOut[17]), .D(n22388), 
         .Z(intgOut0_28__N_735[17])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13563_4_lut_4_lut.init = 16'h00ba;
    LUT4 i2_3_lut_rep_418_4_lut (.A(n6), .B(n21883), .C(n21849), .D(n21848), 
         .Z(n21838)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(174[9:17])
    defparam i2_3_lut_rep_418_4_lut.init = 16'he000;
    LUT4 mux_136_i23_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[22]), 
         .D(backOut1[22]), .Z(n588[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1190_i11_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[10]), 
         .D(speed_set_m3[10]), .Z(n5068)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_136_i7_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[6]), 
         .D(backOut1[6]), .Z(n588[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i28_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[27]), 
         .D(backOut1[27]), .Z(n588[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i28_3_lut_4_lut.init = 16'hfd20;
    AND2 AND2_t64 (.A(subOut[0]), .B(GND_net), .Z(multOut_28__N_1178[0])) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1256[10:66])
    AND2 AND2_t61 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1262[10:66])
    AND2 AND2_t58 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1268[10:66])
    AND2 AND2_t55 (.A(subOut[0]), .B(multIn2[6]), .Z(mult_29s_25s_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1274[10:66])
    AND2 AND2_t52 (.A(subOut[0]), .B(multIn2[6]), .Z(mult_29s_25s_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1280[10:66])
    AND2 AND2_t49 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_5_10)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1286[10:68])
    AND2 AND2_t46 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_6_12)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1292[10:68])
    AND2 AND2_t43 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_7_14)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1298[10:68])
    AND2 AND2_t40 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_8_16)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1304[10:68])
    AND2 AND2_t37 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_9_18)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1310[10:68])
    AND2 AND2_t34 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_10_20)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1316[10:69])
    AND2 AND2_t31 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_11_22)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1322[10:69])
    ND2 ND2_t28 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    ND2 ND2_t27 (.A(subOut[1]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_25)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    ND2 ND2_t26 (.A(subOut[2]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    ND2 ND2_t25 (.A(subOut[3]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_27)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    ND2 ND2_t24 (.A(subOut[4]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 mux_136_i27_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[26]), 
         .D(backOut1[26]), .Z(n588[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i27_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_17_rep_2_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[0]), .B1(subIn2[0]), .C1(GND_net), 
          .D1(GND_net), .COUT(n18754), .S1(n4204));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_1.INIT0 = 16'h0000;
    defparam sub_17_rep_2_add_2_1.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_1.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_1.INJECT1_1 = "NO";
    FADD2B mult_29s_25s_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_12 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_14 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_16 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_18 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_20 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_22 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_0_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_0_2), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_1_2), .CI(GND_net), .COUT(co_mult_29s_25s_0_0_1), 
           .S1(multOut_28__N_1178[2])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_2 (.A0(mult_29s_25s_0_pp_0_3), .A1(mult_29s_25s_0_pp_0_4), 
           .B0(mult_29s_25s_0_pp_1_3), .B1(mult_29s_25s_0_pp_1_4), .CI(co_mult_29s_25s_0_0_1), 
           .COUT(co_mult_29s_25s_0_0_2), .S0(multOut_28__N_1178[3]), .S1(s_mult_29s_25s_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_3 (.A0(mult_29s_25s_0_pp_0_5), .A1(mult_29s_25s_0_pp_0_6), 
           .B0(mult_29s_25s_0_pp_1_5), .B1(mult_29s_25s_0_pp_1_6), .CI(co_mult_29s_25s_0_0_2), 
           .COUT(co_mult_29s_25s_0_0_3), .S0(s_mult_29s_25s_0_0_5), .S1(s_mult_29s_25s_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_4 (.A0(mult_29s_25s_0_pp_0_7), .A1(mult_29s_25s_0_pp_0_8), 
           .B0(mult_29s_25s_0_pp_1_7), .B1(mult_29s_25s_0_pp_1_8), .CI(co_mult_29s_25s_0_0_3), 
           .COUT(co_mult_29s_25s_0_0_4), .S0(s_mult_29s_25s_0_0_7), .S1(s_mult_29s_25s_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_5 (.A0(mult_29s_25s_0_pp_0_9), .A1(mult_29s_25s_0_pp_0_10), 
           .B0(mult_29s_25s_0_pp_1_9), .B1(mult_29s_25s_0_pp_1_10), .CI(co_mult_29s_25s_0_0_4), 
           .COUT(co_mult_29s_25s_0_0_5), .S0(s_mult_29s_25s_0_0_9), .S1(s_mult_29s_25s_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_6 (.A0(mult_29s_25s_0_pp_0_11), .A1(mult_29s_25s_0_pp_0_12), 
           .B0(mult_29s_25s_0_pp_1_11), .B1(mult_29s_25s_0_pp_1_12), .CI(co_mult_29s_25s_0_0_5), 
           .COUT(co_mult_29s_25s_0_0_6), .S0(s_mult_29s_25s_0_0_11), .S1(s_mult_29s_25s_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_7 (.A0(mult_29s_25s_0_pp_0_13), .A1(mult_29s_25s_0_pp_0_14), 
           .B0(mult_29s_25s_0_pp_1_13), .B1(mult_29s_25s_0_pp_1_14), .CI(co_mult_29s_25s_0_0_6), 
           .COUT(co_mult_29s_25s_0_0_7), .S0(s_mult_29s_25s_0_0_13), .S1(s_mult_29s_25s_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_8 (.A0(mult_29s_25s_0_pp_0_15), .A1(mult_29s_25s_0_pp_0_16), 
           .B0(mult_29s_25s_0_pp_1_15), .B1(mult_29s_25s_0_pp_1_16), .CI(co_mult_29s_25s_0_0_7), 
           .COUT(co_mult_29s_25s_0_0_8), .S0(s_mult_29s_25s_0_0_15), .S1(s_mult_29s_25s_0_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_9 (.A0(mult_29s_25s_0_pp_0_17), .A1(mult_29s_25s_0_pp_0_18), 
           .B0(mult_29s_25s_0_pp_1_17), .B1(mult_29s_25s_0_pp_1_18), .CI(co_mult_29s_25s_0_0_8), 
           .COUT(co_mult_29s_25s_0_0_9), .S0(s_mult_29s_25s_0_0_17), .S1(s_mult_29s_25s_0_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_10 (.A0(mult_29s_25s_0_pp_0_19), .A1(mult_29s_25s_0_pp_0_20), 
           .B0(mult_29s_25s_0_pp_1_19), .B1(mult_29s_25s_0_pp_1_20), .CI(co_mult_29s_25s_0_0_9), 
           .COUT(co_mult_29s_25s_0_0_10), .S0(s_mult_29s_25s_0_0_19), .S1(s_mult_29s_25s_0_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_11 (.A0(mult_29s_25s_0_pp_0_21), .A1(mult_29s_25s_0_pp_0_22), 
           .B0(mult_29s_25s_0_pp_1_21), .B1(mult_29s_25s_0_pp_1_22), .CI(co_mult_29s_25s_0_0_10), 
           .COUT(co_mult_29s_25s_0_0_11), .S0(s_mult_29s_25s_0_0_21), .S1(s_mult_29s_25s_0_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_12 (.A0(mult_29s_25s_0_pp_0_23), .A1(mult_29s_25s_0_pp_0_24), 
           .B0(mult_29s_25s_0_pp_1_23), .B1(mult_29s_25s_0_pp_1_24), .CI(co_mult_29s_25s_0_0_11), 
           .COUT(co_mult_29s_25s_0_0_12), .S0(s_mult_29s_25s_0_0_23), .S1(s_mult_29s_25s_0_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_13 (.A0(mult_29s_25s_0_pp_0_25), .A1(mult_29s_25s_0_pp_0_26), 
           .B0(mult_29s_25s_0_pp_1_25), .B1(mult_29s_25s_0_pp_1_26), .CI(co_mult_29s_25s_0_0_12), 
           .COUT(co_mult_29s_25s_0_0_13), .S0(s_mult_29s_25s_0_0_25), .S1(s_mult_29s_25s_0_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_14 (.A0(mult_29s_25s_0_pp_0_27), .A1(mult_29s_25s_0_pp_0_28), 
           .B0(mult_29s_25s_0_pp_1_27), .B1(mult_29s_25s_0_pp_1_28), .CI(co_mult_29s_25s_0_0_13), 
           .S0(s_mult_29s_25s_0_0_27), .S1(s_mult_29s_25s_0_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_1_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_2_6), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_3_6), .CI(GND_net), .COUT(co_mult_29s_25s_0_1_1), 
           .S1(s_mult_29s_25s_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_2 (.A0(mult_29s_25s_0_pp_2_7), .A1(mult_29s_25s_0_pp_2_8), 
           .B0(mult_29s_25s_0_pp_3_7), .B1(mult_29s_25s_0_pp_3_8), .CI(co_mult_29s_25s_0_1_1), 
           .COUT(co_mult_29s_25s_0_1_2), .S0(s_mult_29s_25s_0_1_7), .S1(s_mult_29s_25s_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_3 (.A0(mult_29s_25s_0_pp_2_9), .A1(mult_29s_25s_0_pp_2_10), 
           .B0(mult_29s_25s_0_pp_3_9), .B1(mult_29s_25s_0_pp_3_10), .CI(co_mult_29s_25s_0_1_2), 
           .COUT(co_mult_29s_25s_0_1_3), .S0(s_mult_29s_25s_0_1_9), .S1(s_mult_29s_25s_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_4 (.A0(mult_29s_25s_0_pp_2_11), .A1(mult_29s_25s_0_pp_2_12), 
           .B0(mult_29s_25s_0_pp_3_11), .B1(mult_29s_25s_0_pp_3_12), .CI(co_mult_29s_25s_0_1_3), 
           .COUT(co_mult_29s_25s_0_1_4), .S0(s_mult_29s_25s_0_1_11), .S1(s_mult_29s_25s_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_5 (.A0(mult_29s_25s_0_pp_2_13), .A1(mult_29s_25s_0_pp_2_14), 
           .B0(mult_29s_25s_0_pp_3_13), .B1(mult_29s_25s_0_pp_3_14), .CI(co_mult_29s_25s_0_1_4), 
           .COUT(co_mult_29s_25s_0_1_5), .S0(s_mult_29s_25s_0_1_13), .S1(s_mult_29s_25s_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_6 (.A0(mult_29s_25s_0_pp_2_15), .A1(mult_29s_25s_0_pp_2_16), 
           .B0(mult_29s_25s_0_pp_3_15), .B1(mult_29s_25s_0_pp_3_16), .CI(co_mult_29s_25s_0_1_5), 
           .COUT(co_mult_29s_25s_0_1_6), .S0(s_mult_29s_25s_0_1_15), .S1(s_mult_29s_25s_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_7 (.A0(mult_29s_25s_0_pp_2_17), .A1(mult_29s_25s_0_pp_2_18), 
           .B0(mult_29s_25s_0_pp_3_17), .B1(mult_29s_25s_0_pp_3_18), .CI(co_mult_29s_25s_0_1_6), 
           .COUT(co_mult_29s_25s_0_1_7), .S0(s_mult_29s_25s_0_1_17), .S1(s_mult_29s_25s_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_8 (.A0(mult_29s_25s_0_pp_2_19), .A1(mult_29s_25s_0_pp_2_20), 
           .B0(mult_29s_25s_0_pp_3_19), .B1(mult_29s_25s_0_pp_3_20), .CI(co_mult_29s_25s_0_1_7), 
           .COUT(co_mult_29s_25s_0_1_8), .S0(s_mult_29s_25s_0_1_19), .S1(s_mult_29s_25s_0_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_9 (.A0(mult_29s_25s_0_pp_2_21), .A1(mult_29s_25s_0_pp_2_22), 
           .B0(mult_29s_25s_0_pp_3_21), .B1(mult_29s_25s_0_pp_3_22), .CI(co_mult_29s_25s_0_1_8), 
           .COUT(co_mult_29s_25s_0_1_9), .S0(s_mult_29s_25s_0_1_21), .S1(s_mult_29s_25s_0_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_10 (.A0(mult_29s_25s_0_pp_2_23), .A1(mult_29s_25s_0_pp_2_24), 
           .B0(mult_29s_25s_0_pp_3_23), .B1(mult_29s_25s_0_pp_3_24), .CI(co_mult_29s_25s_0_1_9), 
           .COUT(co_mult_29s_25s_0_1_10), .S0(s_mult_29s_25s_0_1_23), .S1(s_mult_29s_25s_0_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_11 (.A0(mult_29s_25s_0_pp_2_25), .A1(mult_29s_25s_0_pp_2_26), 
           .B0(mult_29s_25s_0_pp_3_25), .B1(mult_29s_25s_0_pp_3_26), .CI(co_mult_29s_25s_0_1_10), 
           .COUT(co_mult_29s_25s_0_1_11), .S0(s_mult_29s_25s_0_1_25), .S1(s_mult_29s_25s_0_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_12 (.A0(mult_29s_25s_0_pp_2_27), .A1(mult_29s_25s_0_pp_2_28), 
           .B0(mult_29s_25s_0_pp_3_27), .B1(mult_29s_25s_0_pp_3_28), .CI(co_mult_29s_25s_0_1_11), 
           .S0(s_mult_29s_25s_0_1_27), .S1(s_mult_29s_25s_0_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 mux_136_i26_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[25]), 
         .D(backOut1[25]), .Z(n588[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i26_3_lut_4_lut.init = 16'hfd20;
    FADD2B Cadd_mult_29s_25s_0_2_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_4_10), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_5_10), .CI(GND_net), .COUT(co_mult_29s_25s_0_2_1), 
           .S1(s_mult_29s_25s_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_2 (.A0(mult_29s_25s_0_pp_4_11), .A1(mult_29s_25s_0_pp_4_12), 
           .B0(mult_29s_25s_0_pp_5_11), .B1(mult_29s_25s_0_pp_5_12), .CI(co_mult_29s_25s_0_2_1), 
           .COUT(co_mult_29s_25s_0_2_2), .S0(s_mult_29s_25s_0_2_11), .S1(s_mult_29s_25s_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_3 (.A0(mult_29s_25s_0_pp_4_13), .A1(mult_29s_25s_0_pp_4_14), 
           .B0(mult_29s_25s_0_pp_5_13), .B1(mult_29s_25s_0_pp_5_14), .CI(co_mult_29s_25s_0_2_2), 
           .COUT(co_mult_29s_25s_0_2_3), .S0(s_mult_29s_25s_0_2_13), .S1(s_mult_29s_25s_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_4 (.A0(mult_29s_25s_0_pp_4_15), .A1(mult_29s_25s_0_pp_4_16), 
           .B0(mult_29s_25s_0_pp_5_15), .B1(mult_29s_25s_0_pp_5_16), .CI(co_mult_29s_25s_0_2_3), 
           .COUT(co_mult_29s_25s_0_2_4), .S0(s_mult_29s_25s_0_2_15), .S1(s_mult_29s_25s_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_5 (.A0(mult_29s_25s_0_pp_4_17), .A1(mult_29s_25s_0_pp_4_18), 
           .B0(mult_29s_25s_0_pp_5_17), .B1(mult_29s_25s_0_pp_5_18), .CI(co_mult_29s_25s_0_2_4), 
           .COUT(co_mult_29s_25s_0_2_5), .S0(s_mult_29s_25s_0_2_17), .S1(s_mult_29s_25s_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_6 (.A0(mult_29s_25s_0_pp_4_19), .A1(mult_29s_25s_0_pp_4_20), 
           .B0(mult_29s_25s_0_pp_5_19), .B1(mult_29s_25s_0_pp_5_20), .CI(co_mult_29s_25s_0_2_5), 
           .COUT(co_mult_29s_25s_0_2_6), .S0(s_mult_29s_25s_0_2_19), .S1(s_mult_29s_25s_0_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_7 (.A0(mult_29s_25s_0_pp_4_21), .A1(mult_29s_25s_0_pp_4_22), 
           .B0(mult_29s_25s_0_pp_5_21), .B1(mult_29s_25s_0_pp_5_22), .CI(co_mult_29s_25s_0_2_6), 
           .COUT(co_mult_29s_25s_0_2_7), .S0(s_mult_29s_25s_0_2_21), .S1(s_mult_29s_25s_0_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_8 (.A0(mult_29s_25s_0_pp_4_23), .A1(mult_29s_25s_0_pp_4_24), 
           .B0(mult_29s_25s_0_pp_5_23), .B1(mult_29s_25s_0_pp_5_24), .CI(co_mult_29s_25s_0_2_7), 
           .COUT(co_mult_29s_25s_0_2_8), .S0(s_mult_29s_25s_0_2_23), .S1(s_mult_29s_25s_0_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_9 (.A0(mult_29s_25s_0_pp_4_25), .A1(mult_29s_25s_0_pp_4_26), 
           .B0(mult_29s_25s_0_pp_5_25), .B1(mult_29s_25s_0_pp_5_26), .CI(co_mult_29s_25s_0_2_8), 
           .COUT(co_mult_29s_25s_0_2_9), .S0(s_mult_29s_25s_0_2_25), .S1(s_mult_29s_25s_0_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_10 (.A0(mult_29s_25s_0_pp_4_27), .A1(mult_29s_25s_0_pp_4_28), 
           .B0(mult_29s_25s_0_pp_5_27), .B1(mult_29s_25s_0_pp_5_28), .CI(co_mult_29s_25s_0_2_9), 
           .S0(s_mult_29s_25s_0_2_27), .S1(s_mult_29s_25s_0_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_3_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_6_14), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_7_14), .CI(GND_net), .COUT(co_mult_29s_25s_0_3_1), 
           .S1(s_mult_29s_25s_0_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_2 (.A0(mult_29s_25s_0_pp_6_15), .A1(mult_29s_25s_0_pp_6_16), 
           .B0(mult_29s_25s_0_pp_7_15), .B1(mult_29s_25s_0_pp_7_16), .CI(co_mult_29s_25s_0_3_1), 
           .COUT(co_mult_29s_25s_0_3_2), .S0(s_mult_29s_25s_0_3_15), .S1(s_mult_29s_25s_0_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_3 (.A0(mult_29s_25s_0_pp_6_17), .A1(mult_29s_25s_0_pp_6_18), 
           .B0(mult_29s_25s_0_pp_7_17), .B1(mult_29s_25s_0_pp_7_18), .CI(co_mult_29s_25s_0_3_2), 
           .COUT(co_mult_29s_25s_0_3_3), .S0(s_mult_29s_25s_0_3_17), .S1(s_mult_29s_25s_0_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_4 (.A0(mult_29s_25s_0_pp_6_19), .A1(mult_29s_25s_0_pp_6_20), 
           .B0(mult_29s_25s_0_pp_7_19), .B1(mult_29s_25s_0_pp_7_20), .CI(co_mult_29s_25s_0_3_3), 
           .COUT(co_mult_29s_25s_0_3_4), .S0(s_mult_29s_25s_0_3_19), .S1(s_mult_29s_25s_0_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_5 (.A0(mult_29s_25s_0_pp_6_21), .A1(mult_29s_25s_0_pp_6_22), 
           .B0(mult_29s_25s_0_pp_7_21), .B1(mult_29s_25s_0_pp_7_22), .CI(co_mult_29s_25s_0_3_4), 
           .COUT(co_mult_29s_25s_0_3_5), .S0(s_mult_29s_25s_0_3_21), .S1(s_mult_29s_25s_0_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_6 (.A0(mult_29s_25s_0_pp_6_23), .A1(mult_29s_25s_0_pp_6_24), 
           .B0(mult_29s_25s_0_pp_7_23), .B1(mult_29s_25s_0_pp_7_24), .CI(co_mult_29s_25s_0_3_5), 
           .COUT(co_mult_29s_25s_0_3_6), .S0(s_mult_29s_25s_0_3_23), .S1(s_mult_29s_25s_0_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_7 (.A0(mult_29s_25s_0_pp_6_25), .A1(mult_29s_25s_0_pp_6_26), 
           .B0(mult_29s_25s_0_pp_7_25), .B1(mult_29s_25s_0_pp_7_26), .CI(co_mult_29s_25s_0_3_6), 
           .COUT(co_mult_29s_25s_0_3_7), .S0(s_mult_29s_25s_0_3_25), .S1(s_mult_29s_25s_0_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_8 (.A0(mult_29s_25s_0_pp_6_27), .A1(mult_29s_25s_0_pp_6_28), 
           .B0(mult_29s_25s_0_pp_7_27), .B1(mult_29s_25s_0_pp_7_28), .CI(co_mult_29s_25s_0_3_7), 
           .S0(s_mult_29s_25s_0_3_27), .S1(s_mult_29s_25s_0_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 i29_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[5]), .D(backOut1[5]), 
         .Z(n10)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam i29_3_lut_4_lut.init = 16'hfd20;
    FADD2B Cadd_mult_29s_25s_0_4_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_8_18), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_9_18), .CI(GND_net), .COUT(co_mult_29s_25s_0_4_1), 
           .S1(s_mult_29s_25s_0_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_2 (.A0(mult_29s_25s_0_pp_8_19), .A1(mult_29s_25s_0_pp_8_20), 
           .B0(mult_29s_25s_0_pp_9_19), .B1(mult_29s_25s_0_pp_9_20), .CI(co_mult_29s_25s_0_4_1), 
           .COUT(co_mult_29s_25s_0_4_2), .S0(s_mult_29s_25s_0_4_19), .S1(s_mult_29s_25s_0_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_3 (.A0(mult_29s_25s_0_pp_8_21), .A1(mult_29s_25s_0_pp_8_22), 
           .B0(mult_29s_25s_0_pp_9_21), .B1(mult_29s_25s_0_pp_9_22), .CI(co_mult_29s_25s_0_4_2), 
           .COUT(co_mult_29s_25s_0_4_3), .S0(s_mult_29s_25s_0_4_21), .S1(s_mult_29s_25s_0_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_4 (.A0(mult_29s_25s_0_pp_8_23), .A1(mult_29s_25s_0_pp_8_24), 
           .B0(mult_29s_25s_0_pp_9_23), .B1(mult_29s_25s_0_pp_9_24), .CI(co_mult_29s_25s_0_4_3), 
           .COUT(co_mult_29s_25s_0_4_4), .S0(s_mult_29s_25s_0_4_23), .S1(s_mult_29s_25s_0_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_5 (.A0(mult_29s_25s_0_pp_8_25), .A1(mult_29s_25s_0_pp_8_26), 
           .B0(mult_29s_25s_0_pp_9_25), .B1(mult_29s_25s_0_pp_9_26), .CI(co_mult_29s_25s_0_4_4), 
           .COUT(co_mult_29s_25s_0_4_5), .S0(s_mult_29s_25s_0_4_25), .S1(s_mult_29s_25s_0_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_6 (.A0(mult_29s_25s_0_pp_8_27), .A1(mult_29s_25s_0_pp_8_28), 
           .B0(mult_29s_25s_0_pp_9_27), .B1(mult_29s_25s_0_pp_9_28), .CI(co_mult_29s_25s_0_4_5), 
           .S0(s_mult_29s_25s_0_4_27), .S1(s_mult_29s_25s_0_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_5_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_10_22), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_11_22), .CI(GND_net), .COUT(co_mult_29s_25s_0_5_1), 
           .S1(s_mult_29s_25s_0_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_2 (.A0(mult_29s_25s_0_pp_10_23), .A1(mult_29s_25s_0_pp_10_24), 
           .B0(mult_29s_25s_0_pp_11_23), .B1(mult_29s_25s_0_pp_11_24), .CI(co_mult_29s_25s_0_5_1), 
           .COUT(co_mult_29s_25s_0_5_2), .S0(s_mult_29s_25s_0_5_23), .S1(s_mult_29s_25s_0_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_3 (.A0(mult_29s_25s_0_pp_10_25), .A1(mult_29s_25s_0_pp_10_26), 
           .B0(mult_29s_25s_0_pp_11_25), .B1(mult_29s_25s_0_pp_11_26), .CI(co_mult_29s_25s_0_5_2), 
           .COUT(co_mult_29s_25s_0_5_3), .S0(s_mult_29s_25s_0_5_25), .S1(s_mult_29s_25s_0_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_4 (.A0(mult_29s_25s_0_pp_10_27), .A1(mult_29s_25s_0_pp_10_28), 
           .B0(mult_29s_25s_0_pp_11_27), .B1(mult_29s_25s_0_pp_11_28), .CI(co_mult_29s_25s_0_5_3), 
           .S0(s_mult_29s_25s_0_5_27), .S1(s_mult_29s_25s_0_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 i29_3_lut_4_lut_adj_39 (.A(n21892), .B(n21868), .C(backOut0[1]), 
         .D(backOut1[1]), .Z(n10_adj_1)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam i29_3_lut_4_lut_adj_39.init = 16'hfd20;
    FADD2B Cadd_mult_29s_25s_0_6_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_12_24), 
           .B0(GND_net), .B1(VCC_net), .CI(GND_net), .COUT(co_mult_29s_25s_0_6_1), 
           .S1(s_mult_29s_25s_0_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_2 (.A0(mult_29s_25s_0_pp_12_25), .A1(mult_29s_25s_0_pp_12_26), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_1), .COUT(co_mult_29s_25s_0_6_2), 
           .S0(s_mult_29s_25s_0_6_25), .S1(s_mult_29s_25s_0_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_3 (.A0(mult_29s_25s_0_pp_12_27), .A1(mult_29s_25s_0_pp_12_28), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_2), .S0(s_mult_29s_25s_0_6_27), 
           .S1(s_mult_29s_25s_0_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 i50_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[0]), .D(backOut1[0]), 
         .Z(n32)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam i50_3_lut_4_lut.init = 16'hfd20;
    FADD2B Cadd_mult_29s_25s_0_7_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_0_4), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_2_4), .CI(GND_net), .COUT(co_mult_29s_25s_0_7_1), 
           .S1(multOut_28__N_1178[4])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_2 (.A0(s_mult_29s_25s_0_0_5), .A1(s_mult_29s_25s_0_0_6), 
           .B0(mult_29s_25s_0_pp_2_5), .B1(s_mult_29s_25s_0_1_6), .CI(co_mult_29s_25s_0_7_1), 
           .COUT(co_mult_29s_25s_0_7_2), .S0(multOut_28__N_1178[5]), .S1(multOut_28__N_1178[6])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_3 (.A0(s_mult_29s_25s_0_0_7), .A1(s_mult_29s_25s_0_0_8), 
           .B0(s_mult_29s_25s_0_1_7), .B1(s_mult_29s_25s_0_1_8), .CI(co_mult_29s_25s_0_7_2), 
           .COUT(co_mult_29s_25s_0_7_3), .S0(multOut_28__N_1178[7]), .S1(s_mult_29s_25s_0_7_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_4 (.A0(s_mult_29s_25s_0_0_9), .A1(s_mult_29s_25s_0_0_10), 
           .B0(s_mult_29s_25s_0_1_9), .B1(s_mult_29s_25s_0_1_10), .CI(co_mult_29s_25s_0_7_3), 
           .COUT(co_mult_29s_25s_0_7_4), .S0(s_mult_29s_25s_0_7_9), .S1(s_mult_29s_25s_0_7_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_5 (.A0(s_mult_29s_25s_0_0_11), .A1(s_mult_29s_25s_0_0_12), 
           .B0(s_mult_29s_25s_0_1_11), .B1(s_mult_29s_25s_0_1_12), .CI(co_mult_29s_25s_0_7_4), 
           .COUT(co_mult_29s_25s_0_7_5), .S0(s_mult_29s_25s_0_7_11), .S1(s_mult_29s_25s_0_7_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_6 (.A0(s_mult_29s_25s_0_0_13), .A1(s_mult_29s_25s_0_0_14), 
           .B0(s_mult_29s_25s_0_1_13), .B1(s_mult_29s_25s_0_1_14), .CI(co_mult_29s_25s_0_7_5), 
           .COUT(co_mult_29s_25s_0_7_6), .S0(s_mult_29s_25s_0_7_13), .S1(s_mult_29s_25s_0_7_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_7 (.A0(s_mult_29s_25s_0_0_15), .A1(s_mult_29s_25s_0_0_16), 
           .B0(s_mult_29s_25s_0_1_15), .B1(s_mult_29s_25s_0_1_16), .CI(co_mult_29s_25s_0_7_6), 
           .COUT(co_mult_29s_25s_0_7_7), .S0(s_mult_29s_25s_0_7_15), .S1(s_mult_29s_25s_0_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_8 (.A0(s_mult_29s_25s_0_0_17), .A1(s_mult_29s_25s_0_0_18), 
           .B0(s_mult_29s_25s_0_1_17), .B1(s_mult_29s_25s_0_1_18), .CI(co_mult_29s_25s_0_7_7), 
           .COUT(co_mult_29s_25s_0_7_8), .S0(s_mult_29s_25s_0_7_17), .S1(s_mult_29s_25s_0_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_9 (.A0(s_mult_29s_25s_0_0_19), .A1(s_mult_29s_25s_0_0_20), 
           .B0(s_mult_29s_25s_0_1_19), .B1(s_mult_29s_25s_0_1_20), .CI(co_mult_29s_25s_0_7_8), 
           .COUT(co_mult_29s_25s_0_7_9), .S0(s_mult_29s_25s_0_7_19), .S1(s_mult_29s_25s_0_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_10 (.A0(s_mult_29s_25s_0_0_21), .A1(s_mult_29s_25s_0_0_22), 
           .B0(s_mult_29s_25s_0_1_21), .B1(s_mult_29s_25s_0_1_22), .CI(co_mult_29s_25s_0_7_9), 
           .COUT(co_mult_29s_25s_0_7_10), .S0(s_mult_29s_25s_0_7_21), .S1(s_mult_29s_25s_0_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_11 (.A0(s_mult_29s_25s_0_0_23), .A1(s_mult_29s_25s_0_0_24), 
           .B0(s_mult_29s_25s_0_1_23), .B1(s_mult_29s_25s_0_1_24), .CI(co_mult_29s_25s_0_7_10), 
           .COUT(co_mult_29s_25s_0_7_11), .S0(s_mult_29s_25s_0_7_23), .S1(s_mult_29s_25s_0_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_12 (.A0(s_mult_29s_25s_0_0_25), .A1(s_mult_29s_25s_0_0_26), 
           .B0(s_mult_29s_25s_0_1_25), .B1(s_mult_29s_25s_0_1_26), .CI(co_mult_29s_25s_0_7_11), 
           .COUT(co_mult_29s_25s_0_7_12), .S0(s_mult_29s_25s_0_7_25), .S1(s_mult_29s_25s_0_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_13 (.A0(s_mult_29s_25s_0_0_27), .A1(s_mult_29s_25s_0_0_28), 
           .B0(s_mult_29s_25s_0_1_27), .B1(s_mult_29s_25s_0_1_28), .CI(co_mult_29s_25s_0_7_12), 
           .S0(s_mult_29s_25s_0_7_27), .S1(s_mult_29s_25s_0_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 mux_1190_i10_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[9]), 
         .D(speed_set_m3[9]), .Z(n5066)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i10_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_mult_29s_25s_0_8_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_2_12), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_6_12), .CI(GND_net), .COUT(co_mult_29s_25s_0_8_1), 
           .S1(s_mult_29s_25s_0_8_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_2 (.A0(s_mult_29s_25s_0_2_13), .A1(s_mult_29s_25s_0_2_14), 
           .B0(mult_29s_25s_0_pp_6_13), .B1(s_mult_29s_25s_0_3_14), .CI(co_mult_29s_25s_0_8_1), 
           .COUT(co_mult_29s_25s_0_8_2), .S0(s_mult_29s_25s_0_8_13), .S1(s_mult_29s_25s_0_8_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_3 (.A0(s_mult_29s_25s_0_2_15), .A1(s_mult_29s_25s_0_2_16), 
           .B0(s_mult_29s_25s_0_3_15), .B1(s_mult_29s_25s_0_3_16), .CI(co_mult_29s_25s_0_8_2), 
           .COUT(co_mult_29s_25s_0_8_3), .S0(s_mult_29s_25s_0_8_15), .S1(s_mult_29s_25s_0_8_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_4 (.A0(s_mult_29s_25s_0_2_17), .A1(s_mult_29s_25s_0_2_18), 
           .B0(s_mult_29s_25s_0_3_17), .B1(s_mult_29s_25s_0_3_18), .CI(co_mult_29s_25s_0_8_3), 
           .COUT(co_mult_29s_25s_0_8_4), .S0(s_mult_29s_25s_0_8_17), .S1(s_mult_29s_25s_0_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_5 (.A0(s_mult_29s_25s_0_2_19), .A1(s_mult_29s_25s_0_2_20), 
           .B0(s_mult_29s_25s_0_3_19), .B1(s_mult_29s_25s_0_3_20), .CI(co_mult_29s_25s_0_8_4), 
           .COUT(co_mult_29s_25s_0_8_5), .S0(s_mult_29s_25s_0_8_19), .S1(s_mult_29s_25s_0_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_6 (.A0(s_mult_29s_25s_0_2_21), .A1(s_mult_29s_25s_0_2_22), 
           .B0(s_mult_29s_25s_0_3_21), .B1(s_mult_29s_25s_0_3_22), .CI(co_mult_29s_25s_0_8_5), 
           .COUT(co_mult_29s_25s_0_8_6), .S0(s_mult_29s_25s_0_8_21), .S1(s_mult_29s_25s_0_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_7 (.A0(s_mult_29s_25s_0_2_23), .A1(s_mult_29s_25s_0_2_24), 
           .B0(s_mult_29s_25s_0_3_23), .B1(s_mult_29s_25s_0_3_24), .CI(co_mult_29s_25s_0_8_6), 
           .COUT(co_mult_29s_25s_0_8_7), .S0(s_mult_29s_25s_0_8_23), .S1(s_mult_29s_25s_0_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_8 (.A0(s_mult_29s_25s_0_2_25), .A1(s_mult_29s_25s_0_2_26), 
           .B0(s_mult_29s_25s_0_3_25), .B1(s_mult_29s_25s_0_3_26), .CI(co_mult_29s_25s_0_8_7), 
           .COUT(co_mult_29s_25s_0_8_8), .S0(s_mult_29s_25s_0_8_25), .S1(s_mult_29s_25s_0_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_9 (.A0(s_mult_29s_25s_0_2_27), .A1(s_mult_29s_25s_0_2_28), 
           .B0(s_mult_29s_25s_0_3_27), .B1(s_mult_29s_25s_0_3_28), .CI(co_mult_29s_25s_0_8_8), 
           .S0(s_mult_29s_25s_0_8_27), .S1(s_mult_29s_25s_0_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 i1_4_lut_4_lut_then_4_lut (.A(ss[2]), .B(ss[3]), .C(ss[0]), .D(ss[1]), 
         .Z(n21926)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_4_lut_then_4_lut.init = 16'hfffe;
    LUT4 mux_1190_i9_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[8]), 
         .D(speed_set_m3[8]), .Z(n5064)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i9_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_mult_29s_25s_0_9_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_4_20), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_10_20), .CI(GND_net), .COUT(co_mult_29s_25s_0_9_1), 
           .S1(s_mult_29s_25s_0_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_2 (.A0(s_mult_29s_25s_0_4_21), .A1(s_mult_29s_25s_0_4_22), 
           .B0(mult_29s_25s_0_pp_10_21), .B1(s_mult_29s_25s_0_5_22), .CI(co_mult_29s_25s_0_9_1), 
           .COUT(co_mult_29s_25s_0_9_2), .S0(s_mult_29s_25s_0_9_21), .S1(s_mult_29s_25s_0_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_3 (.A0(s_mult_29s_25s_0_4_23), .A1(s_mult_29s_25s_0_4_24), 
           .B0(s_mult_29s_25s_0_5_23), .B1(s_mult_29s_25s_0_5_24), .CI(co_mult_29s_25s_0_9_2), 
           .COUT(co_mult_29s_25s_0_9_3), .S0(s_mult_29s_25s_0_9_23), .S1(s_mult_29s_25s_0_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_4 (.A0(s_mult_29s_25s_0_4_25), .A1(s_mult_29s_25s_0_4_26), 
           .B0(s_mult_29s_25s_0_5_25), .B1(s_mult_29s_25s_0_5_26), .CI(co_mult_29s_25s_0_9_3), 
           .COUT(co_mult_29s_25s_0_9_4), .S0(s_mult_29s_25s_0_9_25), .S1(s_mult_29s_25s_0_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_5 (.A0(s_mult_29s_25s_0_4_27), .A1(s_mult_29s_25s_0_4_28), 
           .B0(s_mult_29s_25s_0_5_27), .B1(s_mult_29s_25s_0_5_28), .CI(co_mult_29s_25s_0_9_4), 
           .S0(s_mult_29s_25s_0_9_27), .S1(s_mult_29s_25s_0_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_10_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_7_8), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_4_8), .CI(GND_net), .COUT(co_mult_29s_25s_0_10_1), 
           .S1(multOut_28__N_1178[8])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_2 (.A0(s_mult_29s_25s_0_7_9), .A1(s_mult_29s_25s_0_7_10), 
           .B0(mult_29s_25s_0_pp_4_9), .B1(s_mult_29s_25s_0_2_10), .CI(co_mult_29s_25s_0_10_1), 
           .COUT(co_mult_29s_25s_0_10_2), .S0(multOut_28__N_1178[9]), .S1(multOut_28__N_1178[10])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_3 (.A0(s_mult_29s_25s_0_7_11), .A1(s_mult_29s_25s_0_7_12), 
           .B0(s_mult_29s_25s_0_2_11), .B1(s_mult_29s_25s_0_8_12), .CI(co_mult_29s_25s_0_10_2), 
           .COUT(co_mult_29s_25s_0_10_3), .S0(multOut_28__N_1178[11]), .S1(multOut_28__N_1178[12])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_4 (.A0(s_mult_29s_25s_0_7_13), .A1(s_mult_29s_25s_0_7_14), 
           .B0(s_mult_29s_25s_0_8_13), .B1(s_mult_29s_25s_0_8_14), .CI(co_mult_29s_25s_0_10_3), 
           .COUT(co_mult_29s_25s_0_10_4), .S0(multOut_28__N_1178[13]), .S1(multOut_28__N_1178[14])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_5 (.A0(s_mult_29s_25s_0_7_15), .A1(s_mult_29s_25s_0_7_16), 
           .B0(s_mult_29s_25s_0_8_15), .B1(s_mult_29s_25s_0_8_16), .CI(co_mult_29s_25s_0_10_4), 
           .COUT(co_mult_29s_25s_0_10_5), .S0(multOut_28__N_1178[15]), .S1(s_mult_29s_25s_0_10_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_6 (.A0(s_mult_29s_25s_0_7_17), .A1(s_mult_29s_25s_0_7_18), 
           .B0(s_mult_29s_25s_0_8_17), .B1(s_mult_29s_25s_0_8_18), .CI(co_mult_29s_25s_0_10_5), 
           .COUT(co_mult_29s_25s_0_10_6), .S0(s_mult_29s_25s_0_10_17), .S1(s_mult_29s_25s_0_10_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_7 (.A0(s_mult_29s_25s_0_7_19), .A1(s_mult_29s_25s_0_7_20), 
           .B0(s_mult_29s_25s_0_8_19), .B1(s_mult_29s_25s_0_8_20), .CI(co_mult_29s_25s_0_10_6), 
           .COUT(co_mult_29s_25s_0_10_7), .S0(s_mult_29s_25s_0_10_19), .S1(s_mult_29s_25s_0_10_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_8 (.A0(s_mult_29s_25s_0_7_21), .A1(s_mult_29s_25s_0_7_22), 
           .B0(s_mult_29s_25s_0_8_21), .B1(s_mult_29s_25s_0_8_22), .CI(co_mult_29s_25s_0_10_7), 
           .COUT(co_mult_29s_25s_0_10_8), .S0(s_mult_29s_25s_0_10_21), .S1(s_mult_29s_25s_0_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_9 (.A0(s_mult_29s_25s_0_7_23), .A1(s_mult_29s_25s_0_7_24), 
           .B0(s_mult_29s_25s_0_8_23), .B1(s_mult_29s_25s_0_8_24), .CI(co_mult_29s_25s_0_10_8), 
           .COUT(co_mult_29s_25s_0_10_9), .S0(s_mult_29s_25s_0_10_23), .S1(s_mult_29s_25s_0_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_10 (.A0(s_mult_29s_25s_0_7_25), .A1(s_mult_29s_25s_0_7_26), 
           .B0(s_mult_29s_25s_0_8_25), .B1(s_mult_29s_25s_0_8_26), .CI(co_mult_29s_25s_0_10_9), 
           .COUT(co_mult_29s_25s_0_10_10), .S0(s_mult_29s_25s_0_10_25), 
           .S1(s_mult_29s_25s_0_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_11 (.A0(s_mult_29s_25s_0_7_27), .A1(s_mult_29s_25s_0_7_28), 
           .B0(s_mult_29s_25s_0_8_27), .B1(s_mult_29s_25s_0_8_28), .CI(co_mult_29s_25s_0_10_10), 
           .S0(s_mult_29s_25s_0_10_27), .S1(s_mult_29s_25s_0_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 mux_1190_i8_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[7]), 
         .D(speed_set_m3[7]), .Z(n5062)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1190_i7_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[6]), 
         .D(speed_set_m3[6]), .Z(n5060)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i7_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_mult_29s_25s_0_11_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_9_24), 
           .B0(GND_net), .B1(s_mult_29s_25s_0_6_24), .CI(GND_net), .COUT(co_mult_29s_25s_0_11_1), 
           .S1(s_mult_29s_25s_0_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_2 (.A0(s_mult_29s_25s_0_9_25), .A1(s_mult_29s_25s_0_9_26), 
           .B0(s_mult_29s_25s_0_6_25), .B1(s_mult_29s_25s_0_6_26), .CI(co_mult_29s_25s_0_11_1), 
           .COUT(co_mult_29s_25s_0_11_2), .S0(s_mult_29s_25s_0_11_25), .S1(s_mult_29s_25s_0_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_3 (.A0(s_mult_29s_25s_0_9_27), .A1(s_mult_29s_25s_0_9_28), 
           .B0(s_mult_29s_25s_0_6_27), .B1(s_mult_29s_25s_0_6_28), .CI(co_mult_29s_25s_0_11_2), 
           .S0(s_mult_29s_25s_0_11_27), .S1(s_mult_29s_25s_0_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 i1_2_lut_rep_464_3_lut (.A(ss[0]), .B(ss[2]), .C(ss[1]), .Z(n21884)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_464_3_lut.init = 16'h8080;
    LUT4 i29_3_lut_4_lut_adj_40 (.A(n21892), .B(n21868), .C(backOut0[2]), 
         .D(backOut1[2]), .Z(n10_adj_2)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam i29_3_lut_4_lut_adj_40.init = 16'hfd20;
    FADD2B Cadd_t_mult_29s_25s_0_12_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_10_16), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_8_16), .CI(GND_net), .COUT(co_t_mult_29s_25s_0_12_1), 
           .S1(multOut_28__N_1178[16])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_2 (.A0(s_mult_29s_25s_0_10_17), .A1(s_mult_29s_25s_0_10_18), 
           .B0(mult_29s_25s_0_pp_8_17), .B1(s_mult_29s_25s_0_4_18), .CI(co_t_mult_29s_25s_0_12_1), 
           .COUT(co_t_mult_29s_25s_0_12_2), .S0(multOut_28__N_1178[17]), 
           .S1(multOut_28__N_1178[18])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_3 (.A0(s_mult_29s_25s_0_10_19), .A1(s_mult_29s_25s_0_10_20), 
           .B0(s_mult_29s_25s_0_4_19), .B1(s_mult_29s_25s_0_9_20), .CI(co_t_mult_29s_25s_0_12_2), 
           .COUT(co_t_mult_29s_25s_0_12_3), .S0(multOut_28__N_1178[19]), 
           .S1(multOut_28__N_1178[20])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_4 (.A0(s_mult_29s_25s_0_10_21), .A1(s_mult_29s_25s_0_10_22), 
           .B0(s_mult_29s_25s_0_9_21), .B1(s_mult_29s_25s_0_9_22), .CI(co_t_mult_29s_25s_0_12_3), 
           .COUT(co_t_mult_29s_25s_0_12_4), .S0(multOut_28__N_1178[21]), 
           .S1(multOut_28__N_1178[22])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_5 (.A0(s_mult_29s_25s_0_10_23), .A1(s_mult_29s_25s_0_10_24), 
           .B0(s_mult_29s_25s_0_9_23), .B1(s_mult_29s_25s_0_11_24), .CI(co_t_mult_29s_25s_0_12_4), 
           .COUT(co_t_mult_29s_25s_0_12_5), .S0(multOut_28__N_1178[23]), 
           .S1(multOut_28__N_1178[24])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_6 (.A0(s_mult_29s_25s_0_10_25), .A1(s_mult_29s_25s_0_10_26), 
           .B0(s_mult_29s_25s_0_11_25), .B1(s_mult_29s_25s_0_11_26), .CI(co_t_mult_29s_25s_0_12_5), 
           .COUT(co_t_mult_29s_25s_0_12_6), .S0(multOut_28__N_1178[25]), 
           .S1(multOut_28__N_1178[26])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_7 (.A0(s_mult_29s_25s_0_10_27), .A1(s_mult_29s_25s_0_10_28), 
           .B0(s_mult_29s_25s_0_11_27), .B1(s_mult_29s_25s_0_11_28), .CI(co_t_mult_29s_25s_0_12_6), 
           .S0(multOut_28__N_1178[27]), .S1(multOut_28__N_1178[28])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_0), .CO(mco), .P0(multOut_28__N_1178[1]), 
          .P1(mult_29s_25s_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco), .CO(mco_1), .P0(mult_29s_25s_0_pp_0_3), 
          .P1(mult_29s_25s_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_1), .CO(mco_2), .P0(mult_29s_25s_0_pp_0_5), 
          .P1(mult_29s_25s_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_2), .CO(mco_3), .P0(mult_29s_25s_0_pp_0_7), 
          .P1(mult_29s_25s_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_3), .CO(mco_4), .P0(mult_29s_25s_0_pp_0_9), 
          .P1(mult_29s_25s_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_4), .CO(mco_5), .P0(mult_29s_25s_0_pp_0_11), 
          .P1(mult_29s_25s_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_5), .CO(mco_6), .P0(mult_29s_25s_0_pp_0_13), 
          .P1(mult_29s_25s_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_6), .CO(mco_7), .P0(mult_29s_25s_0_pp_0_15), 
          .P1(mult_29s_25s_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_7), .CO(mco_8), .P0(mult_29s_25s_0_pp_0_17), 
          .P1(mult_29s_25s_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_8), .CO(mco_9), .P0(mult_29s_25s_0_pp_0_19), 
          .P1(mult_29s_25s_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_9), .CO(mco_10), .P0(mult_29s_25s_0_pp_0_21), 
          .P1(mult_29s_25s_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_10), .CO(mco_11), .P0(mult_29s_25s_0_pp_0_23), 
          .P1(mult_29s_25s_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_11), .CO(mco_12), .P0(mult_29s_25s_0_pp_0_25), 
          .P1(mult_29s_25s_0_pp_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_13 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_12), .P0(mult_29s_25s_0_pp_0_27), .P1(mult_29s_25s_0_pp_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_2), .CO(mco_14), 
          .P0(mult_29s_25s_0_pp_1_3), .P1(mult_29s_25s_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_14), .CO(mco_15), .P0(mult_29s_25s_0_pp_1_5), 
          .P1(mult_29s_25s_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_15), .CO(mco_16), .P0(mult_29s_25s_0_pp_1_7), 
          .P1(mult_29s_25s_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_16), .CO(mco_17), .P0(mult_29s_25s_0_pp_1_9), 
          .P1(mult_29s_25s_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_17), .CO(mco_18), .P0(mult_29s_25s_0_pp_1_11), 
          .P1(mult_29s_25s_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_18), .CO(mco_19), .P0(mult_29s_25s_0_pp_1_13), 
          .P1(mult_29s_25s_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_19), .CO(mco_20), .P0(mult_29s_25s_0_pp_1_15), 
          .P1(mult_29s_25s_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_20), .CO(mco_21), .P0(mult_29s_25s_0_pp_1_17), 
          .P1(mult_29s_25s_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_21), .CO(mco_22), .P0(mult_29s_25s_0_pp_1_19), 
          .P1(mult_29s_25s_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_22), .CO(mco_23), .P0(mult_29s_25s_0_pp_1_21), 
          .P1(mult_29s_25s_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_23), .CO(mco_24), .P0(mult_29s_25s_0_pp_1_23), 
          .P1(mult_29s_25s_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_24), .CO(mco_25), .P0(mult_29s_25s_0_pp_1_25), 
          .P1(mult_29s_25s_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_25), .P0(mult_29s_25s_0_pp_1_27), .P1(mult_29s_25s_0_pp_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_4), .CO(mco_28), 
          .P0(mult_29s_25s_0_pp_2_5), .P1(mult_29s_25s_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_28), .CO(mco_29), .P0(mult_29s_25s_0_pp_2_7), 
          .P1(mult_29s_25s_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_29), .CO(mco_30), .P0(mult_29s_25s_0_pp_2_9), 
          .P1(mult_29s_25s_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_30), .CO(mco_31), .P0(mult_29s_25s_0_pp_2_11), 
          .P1(mult_29s_25s_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_31), .CO(mco_32), .P0(mult_29s_25s_0_pp_2_13), 
          .P1(mult_29s_25s_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_32), .CO(mco_33), .P0(mult_29s_25s_0_pp_2_15), 
          .P1(mult_29s_25s_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_33), .CO(mco_34), .P0(mult_29s_25s_0_pp_2_17), 
          .P1(mult_29s_25s_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_34), .CO(mco_35), .P0(mult_29s_25s_0_pp_2_19), 
          .P1(mult_29s_25s_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_35), .CO(mco_36), .P0(mult_29s_25s_0_pp_2_21), 
          .P1(mult_29s_25s_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_36), .CO(mco_37), .P0(mult_29s_25s_0_pp_2_23), 
          .P1(mult_29s_25s_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_37), .CO(mco_38), .P0(mult_29s_25s_0_pp_2_25), 
          .P1(mult_29s_25s_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_38), .P0(mult_29s_25s_0_pp_2_27), .P1(mult_29s_25s_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 i29_3_lut_4_lut_adj_41 (.A(n21892), .B(n21868), .C(backOut0[3]), 
         .D(backOut1[3]), .Z(n10_adj_3)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam i29_3_lut_4_lut_adj_41.init = 16'hfd20;
    MULT2 mult_29s_25s_0_mult_6_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mult_29s_25s_0_cin_lr_6), .CO(mco_42), 
          .P0(mult_29s_25s_0_pp_3_7), .P1(mult_29s_25s_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_42), .CO(mco_43), .P0(mult_29s_25s_0_pp_3_9), 
          .P1(mult_29s_25s_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_43), .CO(mco_44), .P0(mult_29s_25s_0_pp_3_11), 
          .P1(mult_29s_25s_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_44), .CO(mco_45), .P0(mult_29s_25s_0_pp_3_13), 
          .P1(mult_29s_25s_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_45), .CO(mco_46), .P0(mult_29s_25s_0_pp_3_15), 
          .P1(mult_29s_25s_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_46), .CO(mco_47), .P0(mult_29s_25s_0_pp_3_17), 
          .P1(mult_29s_25s_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_47), .CO(mco_48), .P0(mult_29s_25s_0_pp_3_19), 
          .P1(mult_29s_25s_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_48), .CO(mco_49), .P0(mult_29s_25s_0_pp_3_21), 
          .P1(mult_29s_25s_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_49), .CO(mco_50), .P0(mult_29s_25s_0_pp_3_23), 
          .P1(mult_29s_25s_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_50), .CO(mco_51), .P0(mult_29s_25s_0_pp_3_25), 
          .P1(mult_29s_25s_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_51), .P0(mult_29s_25s_0_pp_3_27), .P1(mult_29s_25s_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mult_29s_25s_0_cin_lr_8), .CO(mco_56), 
          .P0(mult_29s_25s_0_pp_4_9), .P1(mult_29s_25s_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_56), .CO(mco_57), .P0(mult_29s_25s_0_pp_4_11), 
          .P1(mult_29s_25s_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_57), .CO(mco_58), .P0(mult_29s_25s_0_pp_4_13), 
          .P1(mult_29s_25s_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_58), .CO(mco_59), .P0(mult_29s_25s_0_pp_4_15), 
          .P1(mult_29s_25s_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_59), .CO(mco_60), .P0(mult_29s_25s_0_pp_4_17), 
          .P1(mult_29s_25s_0_pp_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_60), .CO(mco_61), .P0(mult_29s_25s_0_pp_4_19), 
          .P1(mult_29s_25s_0_pp_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_61), .CO(mco_62), .P0(mult_29s_25s_0_pp_4_21), 
          .P1(mult_29s_25s_0_pp_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_62), .CO(mco_63), .P0(mult_29s_25s_0_pp_4_23), 
          .P1(mult_29s_25s_0_pp_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_63), .CO(mco_64), .P0(mult_29s_25s_0_pp_4_25), 
          .P1(mult_29s_25s_0_pp_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_64), .P0(mult_29s_25s_0_pp_4_27), .P1(mult_29s_25s_0_pp_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_10), .CO(mco_70), .P0(mult_29s_25s_0_pp_5_11), 
          .P1(mult_29s_25s_0_pp_5_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_70), .CO(mco_71), .P0(mult_29s_25s_0_pp_5_13), 
          .P1(mult_29s_25s_0_pp_5_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_71), .CO(mco_72), .P0(mult_29s_25s_0_pp_5_15), 
          .P1(mult_29s_25s_0_pp_5_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_72), .CO(mco_73), .P0(mult_29s_25s_0_pp_5_17), 
          .P1(mult_29s_25s_0_pp_5_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_73), .CO(mco_74), .P0(mult_29s_25s_0_pp_5_19), 
          .P1(mult_29s_25s_0_pp_5_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_74), .CO(mco_75), .P0(mult_29s_25s_0_pp_5_21), 
          .P1(mult_29s_25s_0_pp_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_75), .CO(mco_76), .P0(mult_29s_25s_0_pp_5_23), 
          .P1(mult_29s_25s_0_pp_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_76), .CO(mco_77), .P0(mult_29s_25s_0_pp_5_25), 
          .P1(mult_29s_25s_0_pp_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_77), .P0(mult_29s_25s_0_pp_5_27), .P1(mult_29s_25s_0_pp_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_12), .CO(mco_84), .P0(mult_29s_25s_0_pp_6_13), 
          .P1(mult_29s_25s_0_pp_6_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_84), .CO(mco_85), .P0(mult_29s_25s_0_pp_6_15), 
          .P1(mult_29s_25s_0_pp_6_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_85), .CO(mco_86), .P0(mult_29s_25s_0_pp_6_17), 
          .P1(mult_29s_25s_0_pp_6_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_86), .CO(mco_87), .P0(mult_29s_25s_0_pp_6_19), 
          .P1(mult_29s_25s_0_pp_6_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_87), .CO(mco_88), .P0(mult_29s_25s_0_pp_6_21), 
          .P1(mult_29s_25s_0_pp_6_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_88), .CO(mco_89), .P0(mult_29s_25s_0_pp_6_23), 
          .P1(mult_29s_25s_0_pp_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_89), .CO(mco_90), .P0(mult_29s_25s_0_pp_6_25), 
          .P1(mult_29s_25s_0_pp_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_90), .P0(mult_29s_25s_0_pp_6_27), .P1(mult_29s_25s_0_pp_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 i29_3_lut_4_lut_adj_42 (.A(n21892), .B(n21868), .C(backOut0[4]), 
         .D(backOut1[4]), .Z(n10_adj_4)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam i29_3_lut_4_lut_adj_42.init = 16'hfd20;
    MULT2 mult_29s_25s_0_mult_14_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_14), .CO(mco_98), .P0(mult_29s_25s_0_pp_7_15), 
          .P1(mult_29s_25s_0_pp_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_98), .CO(mco_99), .P0(mult_29s_25s_0_pp_7_17), 
          .P1(mult_29s_25s_0_pp_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_99), .CO(mco_100), .P0(mult_29s_25s_0_pp_7_19), 
          .P1(mult_29s_25s_0_pp_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_100), .CO(mco_101), .P0(mult_29s_25s_0_pp_7_21), 
          .P1(mult_29s_25s_0_pp_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_101), .CO(mco_102), .P0(mult_29s_25s_0_pp_7_23), 
          .P1(mult_29s_25s_0_pp_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_102), .CO(mco_103), .P0(mult_29s_25s_0_pp_7_25), 
          .P1(mult_29s_25s_0_pp_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_103), .P0(mult_29s_25s_0_pp_7_27), .P1(mult_29s_25s_0_pp_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_16), .CO(mco_112), .P0(mult_29s_25s_0_pp_8_17), 
          .P1(mult_29s_25s_0_pp_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_112), .CO(mco_113), .P0(mult_29s_25s_0_pp_8_19), 
          .P1(mult_29s_25s_0_pp_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_113), .CO(mco_114), .P0(mult_29s_25s_0_pp_8_21), 
          .P1(mult_29s_25s_0_pp_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_114), .CO(mco_115), .P0(mult_29s_25s_0_pp_8_23), 
          .P1(mult_29s_25s_0_pp_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_115), .CO(mco_116), .P0(mult_29s_25s_0_pp_8_25), 
          .P1(mult_29s_25s_0_pp_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_116), .P0(mult_29s_25s_0_pp_8_27), .P1(mult_29s_25s_0_pp_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_18), .CO(mco_126), .P0(mult_29s_25s_0_pp_9_19), 
          .P1(mult_29s_25s_0_pp_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_126), .CO(mco_127), .P0(mult_29s_25s_0_pp_9_21), 
          .P1(mult_29s_25s_0_pp_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_127), .CO(mco_128), .P0(mult_29s_25s_0_pp_9_23), 
          .P1(mult_29s_25s_0_pp_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_128), .CO(mco_129), .P0(mult_29s_25s_0_pp_9_25), 
          .P1(mult_29s_25s_0_pp_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_129), .P0(mult_29s_25s_0_pp_9_27), .P1(mult_29s_25s_0_pp_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_20), .CO(mco_140), .P0(mult_29s_25s_0_pp_10_21), 
          .P1(mult_29s_25s_0_pp_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_140), .CO(mco_141), .P0(mult_29s_25s_0_pp_10_23), 
          .P1(mult_29s_25s_0_pp_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_141), .CO(mco_142), .P0(mult_29s_25s_0_pp_10_25), 
          .P1(mult_29s_25s_0_pp_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_142), .P0(mult_29s_25s_0_pp_10_27), .P1(mult_29s_25s_0_pp_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 mux_136_i24_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[23]), 
         .D(backOut1[23]), .Z(n588[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i24_3_lut_4_lut.init = 16'hfd20;
    MULT2 mult_29s_25s_0_mult_22_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_22), .CO(mco_154), .P0(mult_29s_25s_0_pp_11_23), 
          .P1(mult_29s_25s_0_pp_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_154), .CO(mco_155), .P0(mult_29s_25s_0_pp_11_25), 
          .P1(mult_29s_25s_0_pp_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_155), .P0(mult_29s_25s_0_pp_11_27), .P1(mult_29s_25s_0_pp_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 mux_136_i29_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[28]), 
         .D(backOut1[28]), .Z(n588[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1190_i6_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[5]), 
         .D(speed_set_m3[5]), .Z(n5058)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_136_i20_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[19]), 
         .D(backOut1[19]), .Z(n588[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i20_3_lut_4_lut.init = 16'hfd20;
    FADD2B mult_29s_25s_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(229[14:21])
    LUT4 mux_136_i21_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[20]), 
         .D(backOut1[20]), .Z(n588[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_adj_43 (.A(n920), .B(n3636), .C(addOut[4]), 
         .D(n22388), .Z(intgOut0_28__N_735[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_43.init = 16'h0010;
    LUT4 mux_136_i15_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[14]), 
         .D(backOut1[14]), .Z(n588[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i22_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[21]), 
         .D(backOut1[21]), .Z(n588[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i16_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[15]), 
         .D(backOut1[15]), .Z(n588[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 i7_4_lut (.A(Out0[3]), .B(n14_adj_1824), .C(n10_adj_1825), .D(Out0[4]), 
         .Z(n19130)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(ss[3]), .B(n20184), .C(n22388), .D(n21884), .Z(clk_N_683_enable_40)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hc4c0;
    LUT4 mux_136_i9_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[8]), 
         .D(backOut1[8]), .Z(n588[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i17_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[16]), 
         .D(backOut1[16]), .Z(n588[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i6_4_lut (.A(Out0[11]), .B(Out0[7]), .C(Out0[2]), .D(Out0[10]), 
         .Z(n14_adj_1824)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(Out0[9]), .B(Out0[1]), .Z(n10_adj_1825)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 mux_136_i18_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[17]), 
         .D(backOut1[17]), .Z(n588[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i10_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[9]), 
         .D(backOut1[9]), .Z(n588[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 i4_4_lut (.A(Out0[5]), .B(Out0[6]), .C(Out0[0]), .D(n6_adj_1826), 
         .Z(n19131)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 mux_136_i8_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[7]), 
         .D(backOut1[7]), .Z(n588[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i14_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[13]), 
         .D(backOut1[13]), .Z(n588[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i19_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[18]), 
         .D(backOut1[18]), .Z(n588[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut (.A(Out0[8]), .B(Out0[12]), .Z(n6_adj_1826)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam i1_2_lut.init = 16'heeee;
    FD1S3AX addOut_2064__i0 (.D(n121[0]), .CK(clk_N_683), .Q(addOut[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i0.GSR = "ENABLED";
    LUT4 mux_136_i25_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[24]), 
         .D(backOut1[24]), .Z(n588[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i11_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[10]), 
         .D(backOut1[10]), .Z(n588[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i12_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[11]), 
         .D(backOut1[11]), .Z(n588[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i13_3_lut_4_lut (.A(n21892), .B(n21868), .C(backOut0[12]), 
         .D(backOut1[12]), .Z(n588[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(173[9:17])
    defparam mux_136_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1190_i5_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[4]), 
         .D(speed_set_m3[4]), .Z(n5056)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13572_4_lut_4_lut (.A(n920), .B(n3636), .C(addOut[18]), .D(n22388), 
         .Z(intgOut1_28__N_766[18])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13572_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_1190_i4_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[3]), 
         .D(speed_set_m3[3]), .Z(n5054)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3_4_lut (.A(n21820), .B(n21824), .C(n21821), .D(n16074), .Z(n16318)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_4_lut_else_4_lut (.A(ss[2]), .B(ss[3]), .C(ss[0]), .D(ss[1]), 
         .Z(n21925)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_4_lut_else_4_lut.init = 16'h0080;
    LUT4 mux_139_i29_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[28]), 
         .D(n648[28]), .Z(n678[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i10_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[9]), 
         .D(n648[9]), .Z(n678[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i10_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_16120_27 (.A0(addOut[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18908), .COUT(n18909));
    defparam add_16120_27.INIT0 = 16'h0aaa;
    defparam add_16120_27.INIT1 = 16'h0aaa;
    defparam add_16120_27.INJECT1_0 = "NO";
    defparam add_16120_27.INJECT1_1 = "NO";
    CCU2D add_183_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[13]), .B1(n19086), .C1(n19087), .D1(Out1[28]), .COUT(n18690), 
          .S1(n1166[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_1.INIT0 = 16'hF000;
    defparam add_183_1.INIT1 = 16'h56aa;
    defparam add_183_1.INJECT1_0 = "NO";
    defparam add_183_1.INJECT1_1 = "NO";
    FD1P3AX backOut0_i0_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_72), 
            .CK(clk_N_683), .Q(backOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i1.GSR = "DISABLED";
    FD1S3AX multOut_i1 (.D(multOut_28__N_1178[1]), .CK(clk_N_683), .Q(multOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i1.GSR = "ENABLED";
    LUT4 mux_139_i23_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[22]), 
         .D(n648[22]), .Z(n678[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_397_3_lut_4_lut (.A(n21892), .B(n21867), .C(n42), 
         .D(n21836), .Z(n21817)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_397_3_lut_4_lut.init = 16'h20f0;
    LUT4 mux_139_i14_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[13]), 
         .D(n648[13]), .Z(n678[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i21_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[20]), 
         .D(n648[20]), .Z(n678[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13573_4_lut_4_lut (.A(n920), .B(n3636), .C(addOut[19]), .D(n22388), 
         .Z(intgOut1_28__N_766[19])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13573_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_1190_i3_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[2]), 
         .D(speed_set_m3[2]), .Z(n5052)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_139_i20_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[19]), 
         .D(n648[19]), .Z(n678[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1190_i2_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[1]), 
         .D(speed_set_m3[1]), .Z(n5050)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_139_i26_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[25]), 
         .D(n648[25]), .Z(n678[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 i39_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[3]), .D(n23), 
         .Z(n21)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i39_3_lut_4_lut.init = 16'hfd20;
    LUT4 i39_3_lut_4_lut_adj_44 (.A(n21892), .B(n21867), .C(intgOut0[4]), 
         .D(n23_adj_1827), .Z(n21_adj_5)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i39_3_lut_4_lut_adj_44.init = 16'hfd20;
    LUT4 i39_3_lut_4_lut_adj_45 (.A(n21892), .B(n21867), .C(intgOut0[2]), 
         .D(n23_adj_1829), .Z(n21_adj_6)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i39_3_lut_4_lut_adj_45.init = 16'hfd20;
    LUT4 i39_3_lut_4_lut_adj_46 (.A(n21892), .B(n21867), .C(intgOut0[1]), 
         .D(n23_adj_1831), .Z(n21_adj_7)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i39_3_lut_4_lut_adj_46.init = 16'hfd20;
    LUT4 mux_139_i25_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[24]), 
         .D(n648[24]), .Z(n678[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i17_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[16]), 
         .D(n648[16]), .Z(n678[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i7_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[6]), 
         .D(n648[6]), .Z(n678[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i8_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[7]), 
         .D(n648[7]), .Z(n678[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i27_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[26]), 
         .D(n648[26]), .Z(n678[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i19_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[18]), 
         .D(n648[18]), .Z(n678[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i9_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[8]), 
         .D(n648[8]), .Z(n678[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13601_2_lut (.A(addOut[28]), .B(n22388), .Z(backOut2_28__N_1474[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13601_2_lut.init = 16'h2222;
    CCU2D add_16120_25 (.A0(addOut[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18907), .COUT(n18908));
    defparam add_16120_25.INIT0 = 16'h0aaa;
    defparam add_16120_25.INIT1 = 16'h0aaa;
    defparam add_16120_25.INJECT1_0 = "NO";
    defparam add_16120_25.INJECT1_1 = "NO";
    LUT4 i2_4_lut_4_lut (.A(n21815), .B(n21821), .C(n7_c), .D(n16074), 
         .Z(n19454)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam i2_4_lut_4_lut.init = 16'h4000;
    LUT4 mux_139_i18_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[17]), 
         .D(n648[17]), .Z(n678[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i18_3_lut_4_lut.init = 16'hfd20;
    FD1S3AX multOut_i2 (.D(multOut_28__N_1178[2]), .CK(clk_N_683), .Q(multOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i2.GSR = "ENABLED";
    FD1S3AX multOut_i3 (.D(multOut_28__N_1178[3]), .CK(clk_N_683), .Q(multOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i3.GSR = "ENABLED";
    FD1S3AX multOut_i4 (.D(multOut_28__N_1178[4]), .CK(clk_N_683), .Q(multOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i4.GSR = "ENABLED";
    FD1S3AX multOut_i5 (.D(multOut_28__N_1178[5]), .CK(clk_N_683), .Q(multOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i5.GSR = "ENABLED";
    FD1S3AX multOut_i6 (.D(multOut_28__N_1178[6]), .CK(clk_N_683), .Q(multOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i6.GSR = "ENABLED";
    FD1S3AX multOut_i7 (.D(multOut_28__N_1178[7]), .CK(clk_N_683), .Q(multOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i7.GSR = "ENABLED";
    FD1S3AX multOut_i8 (.D(multOut_28__N_1178[8]), .CK(clk_N_683), .Q(multOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i8.GSR = "ENABLED";
    FD1S3AX multOut_i9 (.D(multOut_28__N_1178[9]), .CK(clk_N_683), .Q(multOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i9.GSR = "ENABLED";
    FD1S3AX multOut_i10 (.D(multOut_28__N_1178[10]), .CK(clk_N_683), .Q(multOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i10.GSR = "ENABLED";
    FD1S3AX multOut_i11 (.D(multOut_28__N_1178[11]), .CK(clk_N_683), .Q(multOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i11.GSR = "ENABLED";
    FD1S3AX multOut_i12 (.D(multOut_28__N_1178[12]), .CK(clk_N_683), .Q(multOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i12.GSR = "ENABLED";
    FD1S3AX multOut_i13 (.D(multOut_28__N_1178[13]), .CK(clk_N_683), .Q(multOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i13.GSR = "ENABLED";
    FD1S3AX multOut_i14 (.D(multOut_28__N_1178[14]), .CK(clk_N_683), .Q(multOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i14.GSR = "ENABLED";
    FD1S3AX multOut_i15 (.D(multOut_28__N_1178[15]), .CK(clk_N_683), .Q(multOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i15.GSR = "ENABLED";
    FD1S3AX multOut_i16 (.D(multOut_28__N_1178[16]), .CK(clk_N_683), .Q(multOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i16.GSR = "ENABLED";
    FD1S3AX multOut_i17 (.D(multOut_28__N_1178[17]), .CK(clk_N_683), .Q(multOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i17.GSR = "ENABLED";
    FD1S3AX multOut_i18 (.D(multOut_28__N_1178[18]), .CK(clk_N_683), .Q(multOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i18.GSR = "ENABLED";
    FD1S3AX multOut_i19 (.D(multOut_28__N_1178[19]), .CK(clk_N_683), .Q(multOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i19.GSR = "ENABLED";
    FD1S3AX multOut_i20 (.D(multOut_28__N_1178[20]), .CK(clk_N_683), .Q(multOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i20.GSR = "ENABLED";
    FD1S3AX multOut_i21 (.D(multOut_28__N_1178[21]), .CK(clk_N_683), .Q(multOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i21.GSR = "ENABLED";
    FD1S3AX multOut_i22 (.D(multOut_28__N_1178[22]), .CK(clk_N_683), .Q(multOut[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i22.GSR = "ENABLED";
    FD1S3AX multOut_i23 (.D(multOut_28__N_1178[23]), .CK(clk_N_683), .Q(multOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i23.GSR = "ENABLED";
    FD1S3AX multOut_i24 (.D(multOut_28__N_1178[24]), .CK(clk_N_683), .Q(multOut[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i24.GSR = "ENABLED";
    FD1S3AX multOut_i25 (.D(multOut_28__N_1178[25]), .CK(clk_N_683), .Q(multOut[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i25.GSR = "ENABLED";
    FD1S3AX multOut_i26 (.D(multOut_28__N_1178[26]), .CK(clk_N_683), .Q(multOut[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i26.GSR = "ENABLED";
    FD1S3AX multOut_i27 (.D(multOut_28__N_1178[27]), .CK(clk_N_683), .Q(multOut[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i27.GSR = "ENABLED";
    FD1S3AX multOut_i28 (.D(multOut_28__N_1178[28]), .CK(clk_N_683), .Q(multOut[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam multOut_i28.GSR = "ENABLED";
    FD1P3AX intgOut0_i1 (.D(intgOut1_28__N_766[1]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i1.GSR = "ENABLED";
    FD1P3AX intgOut0_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i2.GSR = "ENABLED";
    FD1P3AX intgOut0_i3 (.D(intgOut1_28__N_766[3]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i3.GSR = "ENABLED";
    FD1P3AX intgOut0_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i4.GSR = "ENABLED";
    FD1P3AX intgOut0_i5 (.D(intgOut1_28__N_766[5]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i5.GSR = "ENABLED";
    FD1P3AX intgOut0_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i6.GSR = "ENABLED";
    FD1P3AX intgOut0_i7 (.D(intgOut1_28__N_766[7]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i7.GSR = "ENABLED";
    FD1P3AX intgOut0_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i8.GSR = "ENABLED";
    FD1P3AX intgOut0_i9 (.D(intgOut1_28__N_766[9]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i9.GSR = "ENABLED";
    FD1P3AX intgOut0_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i10.GSR = "ENABLED";
    FD1P3AX intgOut0_i11 (.D(intgOut1_28__N_766[11]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i11.GSR = "ENABLED";
    FD1P3AX intgOut0_i12 (.D(intgOut1_28__N_766[12]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i12.GSR = "ENABLED";
    FD1P3AX intgOut0_i13 (.D(intgOut1_28__N_766[13]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i13.GSR = "ENABLED";
    FD1P3AX intgOut0_i14 (.D(intgOut1_28__N_766[14]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i14.GSR = "ENABLED";
    FD1P3AX intgOut0_i15 (.D(intgOut2_28__N_795[15]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i15.GSR = "ENABLED";
    FD1P3AX intgOut0_i16 (.D(intgOut1_28__N_766[16]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i16.GSR = "ENABLED";
    FD1P3AX intgOut0_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i17.GSR = "ENABLED";
    FD1P3AX intgOut0_i18 (.D(intgOut1_28__N_766[18]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i18.GSR = "ENABLED";
    FD1P3AX intgOut0_i19 (.D(intgOut1_28__N_766[19]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i19.GSR = "ENABLED";
    FD1P3AX intgOut0_i20 (.D(intgOut1_28__N_766[20]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i20.GSR = "ENABLED";
    FD1P3AX intgOut0_i21 (.D(intgOut1_28__N_766[21]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i21.GSR = "ENABLED";
    FD1P3AX intgOut0_i22 (.D(intgOut2_28__N_795[22]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i22.GSR = "ENABLED";
    FD1P3AX intgOut0_i23 (.D(intgOut1_28__N_766[23]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i23.GSR = "ENABLED";
    FD1P3AX intgOut0_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i24.GSR = "ENABLED";
    FD1P3AX intgOut0_i25 (.D(intgOut1_28__N_766[25]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i25.GSR = "ENABLED";
    FD1P3AX intgOut0_i26 (.D(intgOut1_28__N_766[26]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i26.GSR = "ENABLED";
    FD1P3AX intgOut0_i27 (.D(intgOut1_28__N_766[27]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i27.GSR = "ENABLED";
    FD1P3AX intgOut0_i28 (.D(intgOut1_28__N_766[28]), .SP(clk_N_683_enable_100), 
            .CK(clk_N_683), .Q(intgOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut0_i28.GSR = "ENABLED";
    FD1P3AX intgOut1_i1 (.D(intgOut1_28__N_766[1]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i1.GSR = "ENABLED";
    FD1P3AX intgOut1_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i2.GSR = "ENABLED";
    FD1P3AX intgOut1_i3 (.D(intgOut1_28__N_766[3]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i3.GSR = "ENABLED";
    FD1P3AX intgOut1_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i4.GSR = "ENABLED";
    FD1P3AX intgOut1_i5 (.D(intgOut1_28__N_766[5]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i5.GSR = "ENABLED";
    FD1P3AX intgOut1_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i6.GSR = "ENABLED";
    FD1P3AX intgOut1_i7 (.D(intgOut1_28__N_766[7]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i7.GSR = "ENABLED";
    FD1P3AX intgOut1_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i8.GSR = "ENABLED";
    FD1P3AX intgOut1_i9 (.D(intgOut1_28__N_766[9]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i9.GSR = "ENABLED";
    FD1P3AX intgOut1_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i10.GSR = "ENABLED";
    FD1P3AX intgOut1_i11 (.D(intgOut1_28__N_766[11]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i11.GSR = "ENABLED";
    FD1P3AX intgOut1_i12 (.D(intgOut1_28__N_766[12]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i12.GSR = "ENABLED";
    FD1P3AX intgOut1_i13 (.D(intgOut1_28__N_766[13]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i13.GSR = "ENABLED";
    FD1P3AX intgOut1_i14 (.D(intgOut1_28__N_766[14]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i14.GSR = "ENABLED";
    FD1P3AX intgOut1_i15 (.D(intgOut2_28__N_795[15]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i15.GSR = "ENABLED";
    FD1P3AX intgOut1_i16 (.D(intgOut1_28__N_766[16]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i16.GSR = "ENABLED";
    FD1P3AX intgOut1_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i17.GSR = "ENABLED";
    FD1P3AX intgOut1_i18 (.D(intgOut1_28__N_766[18]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i18.GSR = "ENABLED";
    FD1P3AX intgOut1_i19 (.D(intgOut1_28__N_766[19]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i19.GSR = "ENABLED";
    FD1P3AX intgOut1_i20 (.D(intgOut1_28__N_766[20]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i20.GSR = "ENABLED";
    FD1P3AX intgOut1_i21 (.D(intgOut1_28__N_766[21]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i21.GSR = "ENABLED";
    FD1P3AX intgOut1_i22 (.D(intgOut2_28__N_795[22]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i22.GSR = "ENABLED";
    FD1P3AX intgOut1_i23 (.D(intgOut1_28__N_766[23]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i23.GSR = "ENABLED";
    FD1P3AX intgOut1_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i24.GSR = "ENABLED";
    FD1P3AX intgOut1_i25 (.D(intgOut1_28__N_766[25]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i25.GSR = "ENABLED";
    FD1P3AX intgOut1_i26 (.D(intgOut1_28__N_766[26]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i26.GSR = "ENABLED";
    FD1P3AX intgOut1_i27 (.D(intgOut1_28__N_766[27]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i27.GSR = "ENABLED";
    FD1P3AX intgOut1_i28 (.D(intgOut1_28__N_766[28]), .SP(clk_N_683_enable_128), 
            .CK(clk_N_683), .Q(intgOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut1_i28.GSR = "ENABLED";
    FD1P3AX intgOut2_i1 (.D(intgOut1_28__N_766[1]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i1.GSR = "ENABLED";
    FD1P3AX intgOut2_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i2.GSR = "ENABLED";
    FD1P3AX intgOut2_i3 (.D(intgOut1_28__N_766[3]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i3.GSR = "ENABLED";
    FD1P3AX intgOut2_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i4.GSR = "ENABLED";
    FD1P3AX intgOut2_i5 (.D(intgOut1_28__N_766[5]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i5.GSR = "ENABLED";
    FD1P3AX intgOut2_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i6.GSR = "ENABLED";
    FD1P3AX intgOut2_i7 (.D(intgOut1_28__N_766[7]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i7.GSR = "ENABLED";
    FD1P3AX intgOut2_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i8.GSR = "ENABLED";
    FD1P3AX intgOut2_i9 (.D(intgOut1_28__N_766[9]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i9.GSR = "ENABLED";
    FD1P3AX intgOut2_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i10.GSR = "ENABLED";
    FD1P3AX intgOut2_i11 (.D(intgOut1_28__N_766[11]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i11.GSR = "ENABLED";
    FD1P3AX intgOut2_i12 (.D(intgOut1_28__N_766[12]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i12.GSR = "ENABLED";
    FD1P3AX intgOut2_i13 (.D(intgOut1_28__N_766[13]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i13.GSR = "ENABLED";
    FD1P3AX intgOut2_i14 (.D(intgOut1_28__N_766[14]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i14.GSR = "ENABLED";
    FD1P3AX intgOut2_i15 (.D(intgOut2_28__N_795[15]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i15.GSR = "ENABLED";
    FD1P3AX intgOut2_i16 (.D(intgOut1_28__N_766[16]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i16.GSR = "ENABLED";
    FD1P3AX intgOut2_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i17.GSR = "ENABLED";
    FD1P3AX intgOut2_i18 (.D(intgOut1_28__N_766[18]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i18.GSR = "ENABLED";
    FD1P3AX intgOut2_i19 (.D(intgOut1_28__N_766[19]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i19.GSR = "ENABLED";
    FD1P3AX intgOut2_i20 (.D(intgOut1_28__N_766[20]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i20.GSR = "ENABLED";
    FD1P3AX intgOut2_i21 (.D(intgOut1_28__N_766[21]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i21.GSR = "ENABLED";
    FD1P3AX intgOut2_i22 (.D(intgOut2_28__N_795[22]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i22.GSR = "ENABLED";
    FD1P3AX intgOut2_i23 (.D(intgOut1_28__N_766[23]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i23.GSR = "ENABLED";
    FD1P3AX intgOut2_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i24.GSR = "ENABLED";
    FD1P3AX intgOut2_i25 (.D(intgOut1_28__N_766[25]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i25.GSR = "ENABLED";
    FD1P3AX intgOut2_i26 (.D(intgOut1_28__N_766[26]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i26.GSR = "ENABLED";
    FD1P3AX intgOut2_i27 (.D(intgOut1_28__N_766[27]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i27.GSR = "ENABLED";
    FD1P3AX intgOut2_i28 (.D(intgOut1_28__N_766[28]), .SP(clk_N_683_enable_156), 
            .CK(clk_N_683), .Q(intgOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut2_i28.GSR = "ENABLED";
    FD1P3AX intgOut3_i1 (.D(intgOut1_28__N_766[1]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i1.GSR = "ENABLED";
    FD1P3AX intgOut3_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i2.GSR = "ENABLED";
    FD1P3AX intgOut3_i3 (.D(intgOut1_28__N_766[3]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i3.GSR = "ENABLED";
    FD1P3AX intgOut3_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i4.GSR = "ENABLED";
    FD1P3AX intgOut3_i5 (.D(intgOut1_28__N_766[5]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i5.GSR = "ENABLED";
    FD1P3AX intgOut3_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i6.GSR = "ENABLED";
    FD1P3AX intgOut3_i7 (.D(intgOut1_28__N_766[7]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i7.GSR = "ENABLED";
    FD1P3AX intgOut3_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i8.GSR = "ENABLED";
    FD1P3AX intgOut3_i9 (.D(intgOut1_28__N_766[9]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i9.GSR = "ENABLED";
    FD1P3AX intgOut3_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i10.GSR = "ENABLED";
    FD1P3AX intgOut3_i11 (.D(intgOut1_28__N_766[11]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i11.GSR = "ENABLED";
    FD1P3AX intgOut3_i12 (.D(intgOut1_28__N_766[12]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i12.GSR = "ENABLED";
    FD1P3AX intgOut3_i13 (.D(intgOut1_28__N_766[13]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i13.GSR = "ENABLED";
    FD1P3AX intgOut3_i14 (.D(intgOut1_28__N_766[14]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i14.GSR = "ENABLED";
    FD1P3AX intgOut3_i15 (.D(intgOut2_28__N_795[15]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i15.GSR = "ENABLED";
    FD1P3AX intgOut3_i16 (.D(intgOut1_28__N_766[16]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i16.GSR = "ENABLED";
    FD1P3AX intgOut3_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i17.GSR = "ENABLED";
    FD1P3AX intgOut3_i18 (.D(intgOut1_28__N_766[18]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i18.GSR = "ENABLED";
    FD1P3AX intgOut3_i19 (.D(intgOut1_28__N_766[19]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i19.GSR = "ENABLED";
    FD1P3AX intgOut3_i20 (.D(intgOut1_28__N_766[20]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i20.GSR = "ENABLED";
    FD1P3AX intgOut3_i21 (.D(intgOut1_28__N_766[21]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i21.GSR = "ENABLED";
    FD1P3AX intgOut3_i22 (.D(intgOut2_28__N_795[22]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i22.GSR = "ENABLED";
    FD1P3AX intgOut3_i23 (.D(intgOut1_28__N_766[23]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i23.GSR = "ENABLED";
    FD1P3AX intgOut3_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i24.GSR = "ENABLED";
    FD1P3AX intgOut3_i25 (.D(intgOut1_28__N_766[25]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i25.GSR = "ENABLED";
    FD1P3AX intgOut3_i26 (.D(intgOut1_28__N_766[26]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i26.GSR = "ENABLED";
    FD1P3AX intgOut3_i27 (.D(intgOut1_28__N_766[27]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i27.GSR = "ENABLED";
    FD1P3AX intgOut3_i28 (.D(intgOut1_28__N_766[28]), .SP(clk_N_683_enable_184), 
            .CK(clk_N_683), .Q(intgOut3_c[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam intgOut3_i28.GSR = "ENABLED";
    FD1P3AX Out0_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i1.GSR = "ENABLED";
    FD1P3AX Out0_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i2.GSR = "ENABLED";
    FD1P3AX Out0_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i3.GSR = "ENABLED";
    FD1P3AX Out0_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i4.GSR = "ENABLED";
    FD1P3AX Out0_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i5.GSR = "ENABLED";
    FD1P3AX Out0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i6.GSR = "ENABLED";
    FD1P3AX Out0_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_212), .CK(clk_N_683), 
            .Q(Out0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i7.GSR = "ENABLED";
    FD1P3AX Out0_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i8.GSR = "ENABLED";
    FD1P3AX Out0_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i9.GSR = "ENABLED";
    FD1P3AX Out0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i10.GSR = "ENABLED";
    FD1P3AX Out0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i11.GSR = "ENABLED";
    FD1P3AX Out0_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i12.GSR = "ENABLED";
    FD1P3AX Out0_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i13.GSR = "ENABLED";
    FD1P3AX Out0_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i14.GSR = "ENABLED";
    FD1P3AX Out0_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i15.GSR = "ENABLED";
    FD1P3AX Out0_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i16.GSR = "ENABLED";
    FD1P3AX Out0_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i17.GSR = "ENABLED";
    FD1P3AX Out0_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i18.GSR = "ENABLED";
    FD1P3AX Out0_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i19.GSR = "ENABLED";
    FD1P3AX Out0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i20.GSR = "ENABLED";
    FD1P3AX Out0_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i21.GSR = "ENABLED";
    FD1P3AX Out0_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i22.GSR = "ENABLED";
    FD1P3AX Out0_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i23.GSR = "ENABLED";
    FD1P3AX Out0_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i24.GSR = "ENABLED";
    FD1P3AX Out0_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i25.GSR = "ENABLED";
    FD1P3AX Out0_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i26.GSR = "ENABLED";
    FD1P3AX Out0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i27.GSR = "ENABLED";
    FD1P3AX Out0_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_212), 
            .CK(clk_N_683), .Q(Out0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out0_i28.GSR = "ENABLED";
    FD1P3AX Out1_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i1.GSR = "ENABLED";
    FD1P3AX Out1_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i2.GSR = "ENABLED";
    FD1P3AX Out1_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i3.GSR = "ENABLED";
    FD1P3AX Out1_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i4.GSR = "ENABLED";
    FD1P3AX Out1_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i5.GSR = "ENABLED";
    FD1P3AX Out1_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i6.GSR = "ENABLED";
    FD1P3AX Out1_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_240), .CK(clk_N_683), 
            .Q(Out1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i7.GSR = "ENABLED";
    FD1P3AX Out1_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i8.GSR = "ENABLED";
    FD1P3AX Out1_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i9.GSR = "ENABLED";
    FD1P3AX Out1_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i10.GSR = "ENABLED";
    FD1P3AX Out1_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i11.GSR = "ENABLED";
    FD1P3AX Out1_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i12.GSR = "ENABLED";
    FD1P3AX Out1_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i13.GSR = "ENABLED";
    FD1P3AX Out1_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i14.GSR = "ENABLED";
    FD1P3AX Out1_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i15.GSR = "ENABLED";
    FD1P3AX Out1_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i16.GSR = "ENABLED";
    FD1P3AX Out1_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i17.GSR = "ENABLED";
    FD1P3AX Out1_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i18.GSR = "ENABLED";
    FD1P3AX Out1_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i19.GSR = "ENABLED";
    FD1P3AX Out1_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i20.GSR = "ENABLED";
    FD1P3AX Out1_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i21.GSR = "ENABLED";
    FD1P3AX Out1_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i22.GSR = "ENABLED";
    FD1P3AX Out1_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i23.GSR = "ENABLED";
    FD1P3AX Out1_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i24.GSR = "ENABLED";
    FD1P3AX Out1_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i25.GSR = "ENABLED";
    FD1P3AX Out1_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i26.GSR = "ENABLED";
    FD1P3AX Out1_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i27.GSR = "ENABLED";
    FD1P3AX Out1_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_240), 
            .CK(clk_N_683), .Q(Out1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out1_i28.GSR = "ENABLED";
    FD1P3AX Out2_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i1.GSR = "ENABLED";
    FD1P3AX Out2_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i2.GSR = "ENABLED";
    FD1P3AX Out2_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i3.GSR = "ENABLED";
    FD1P3AX Out2_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i4.GSR = "ENABLED";
    FD1P3AX Out2_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i5.GSR = "ENABLED";
    FD1P3AX Out2_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i6.GSR = "ENABLED";
    FD1P3AX Out2_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_268), .CK(clk_N_683), 
            .Q(Out2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i7.GSR = "ENABLED";
    FD1P3AX Out2_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i8.GSR = "ENABLED";
    FD1P3AX Out2_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i9.GSR = "ENABLED";
    FD1P3AX Out2_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i10.GSR = "ENABLED";
    FD1P3AX Out2_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i11.GSR = "ENABLED";
    FD1P3AX Out2_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i12.GSR = "ENABLED";
    FD1P3AX Out2_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i13.GSR = "ENABLED";
    FD1P3AX Out2_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i14.GSR = "ENABLED";
    FD1P3AX Out2_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i15.GSR = "ENABLED";
    FD1P3AX Out2_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i16.GSR = "ENABLED";
    FD1P3AX Out2_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i17.GSR = "ENABLED";
    FD1P3AX Out2_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i18.GSR = "ENABLED";
    FD1P3AX Out2_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i19.GSR = "ENABLED";
    FD1P3AX Out2_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i20.GSR = "ENABLED";
    FD1P3AX Out2_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i21.GSR = "ENABLED";
    FD1P3AX Out2_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i22.GSR = "ENABLED";
    FD1P3AX Out2_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i23.GSR = "ENABLED";
    FD1P3AX Out2_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i24.GSR = "ENABLED";
    FD1P3AX Out2_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i25.GSR = "ENABLED";
    FD1P3AX Out2_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i26.GSR = "ENABLED";
    FD1P3AX Out2_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i27.GSR = "ENABLED";
    FD1P3AX Out2_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_268), 
            .CK(clk_N_683), .Q(Out2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out2_i28.GSR = "ENABLED";
    FD1P3AX Out3_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i1.GSR = "ENABLED";
    FD1P3AX Out3_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i2.GSR = "ENABLED";
    FD1P3AX Out3_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i3.GSR = "ENABLED";
    FD1P3AX Out3_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i4.GSR = "ENABLED";
    FD1P3AX Out3_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i5.GSR = "ENABLED";
    FD1P3AX Out3_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i6.GSR = "ENABLED";
    FD1P3AX Out3_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_296), .CK(clk_N_683), 
            .Q(Out3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i7.GSR = "ENABLED";
    FD1P3AX Out3_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i8.GSR = "ENABLED";
    FD1P3AX Out3_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i9.GSR = "ENABLED";
    FD1P3AX Out3_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i10.GSR = "ENABLED";
    FD1P3AX Out3_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i11.GSR = "ENABLED";
    FD1P3AX Out3_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i12.GSR = "ENABLED";
    FD1P3AX Out3_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i13.GSR = "ENABLED";
    FD1P3AX Out3_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i14.GSR = "ENABLED";
    FD1P3AX Out3_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i15.GSR = "ENABLED";
    FD1P3AX Out3_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i16.GSR = "ENABLED";
    FD1P3AX Out3_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i17.GSR = "ENABLED";
    FD1P3AX Out3_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i18.GSR = "ENABLED";
    FD1P3AX Out3_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i19.GSR = "ENABLED";
    FD1P3AX Out3_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i20.GSR = "ENABLED";
    FD1P3AX Out3_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i21.GSR = "ENABLED";
    FD1P3AX Out3_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i22.GSR = "ENABLED";
    FD1P3AX Out3_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i23.GSR = "ENABLED";
    FD1P3AX Out3_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i24.GSR = "ENABLED";
    FD1P3AX Out3_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i25.GSR = "ENABLED";
    FD1P3AX Out3_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i26.GSR = "ENABLED";
    FD1P3AX Out3_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i27.GSR = "ENABLED";
    FD1P3AX Out3_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_296), 
            .CK(clk_N_683), .Q(Out3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam Out3_i28.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_324), 
            .CK(clk_N_683), .Q(backOut2_c[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i1 (.D(backOut2_28__N_1474[1]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i2 (.D(backOut3_28__N_1503[2]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i3 (.D(backOut2_28__N_1474[3]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i4 (.D(backOut1_28__N_1445[4]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i5 (.D(backOut2_28__N_1474[5]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i7 (.D(Out0_28__N_853[7]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i8 (.D(backOut2_28__N_1474[8]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i9 (.D(backOut2_28__N_1474[9]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i12 (.D(backOut1_28__N_1445[12]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i13 (.D(backOut1_28__N_1445[13]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i14 (.D(backOut2_28__N_1474[14]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i15 (.D(backOut2_28__N_1474[15]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i16 (.D(backOut2_28__N_1474[16]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i17 (.D(backOut3_28__N_1503[17]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i18 (.D(backOut2_28__N_1474[18]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i19 (.D(backOut1_28__N_1445[19]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i21 (.D(backOut2_28__N_1474[21]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i22 (.D(backOut2_28__N_1474[22]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i23 (.D(backOut2_28__N_1474[23]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i24 (.D(backOut3_28__N_1503[24]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i25 (.D(backOut2_28__N_1474[25]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i26 (.D(backOut1_28__N_1445[26]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i28 (.D(backOut2_28__N_1474[28]), .SP(clk_N_683_enable_352), 
            .CK(clk_N_683), .Q(backOut3_c[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i28.GSR = "DISABLED";
    LUT4 i13589_2_lut (.A(addOut[27]), .B(n22388), .Z(backOut1_28__N_1445[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13589_2_lut.init = 16'h2222;
    LUT4 mux_139_i24_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[23]), 
         .D(n648[23]), .Z(n678[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 i39_3_lut_4_lut_adj_47 (.A(n21892), .B(n21867), .C(intgOut0[5]), 
         .D(n23_adj_1833), .Z(n21_adj_8)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i39_3_lut_4_lut_adj_47.init = 16'hfd20;
    LUT4 mux_139_i13_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[12]), 
         .D(n648[12]), .Z(n678[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 i14031_2_lut_rep_400_3_lut_4_lut (.A(n21892), .B(n21867), .C(n42), 
         .D(n21836), .Z(n21820)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C+(D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i14031_2_lut_rep_400_3_lut_4_lut.init = 16'hfdf0;
    LUT4 i48_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[0]), .D(n28), 
         .Z(n30)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam i48_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13588_2_lut (.A(addOut[26]), .B(n22388), .Z(backOut1_28__N_1445[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13588_2_lut.init = 16'h2222;
    LUT4 mux_139_i22_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[21]), 
         .D(n648[21]), .Z(n678[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i22_3_lut_4_lut.init = 16'hfd20;
    FD1S3AX subOut_i1 (.D(\subOut_24__N_1135[1] ), .CK(clk_N_683), .Q(subOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i1.GSR = "ENABLED";
    FD1S3AX subOut_i2 (.D(\subOut_24__N_1135[2] ), .CK(clk_N_683), .Q(subOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i2.GSR = "ENABLED";
    FD1S3AX subOut_i3 (.D(\subOut_24__N_1135[3] ), .CK(clk_N_683), .Q(subOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i3.GSR = "ENABLED";
    FD1S3AX subOut_i4 (.D(\subOut_24__N_1135[4] ), .CK(clk_N_683), .Q(subOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i4.GSR = "ENABLED";
    FD1S3AX subOut_i5 (.D(\subOut_24__N_1135[5] ), .CK(clk_N_683), .Q(subOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i5.GSR = "ENABLED";
    FD1S3AX subOut_i6 (.D(\subOut_24__N_1135[6] ), .CK(clk_N_683), .Q(subOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i6.GSR = "ENABLED";
    FD1S3AX subOut_i7 (.D(\subOut_24__N_1135[7] ), .CK(clk_N_683), .Q(subOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i7.GSR = "ENABLED";
    FD1S3AX subOut_i8 (.D(\subOut_24__N_1135[8] ), .CK(clk_N_683), .Q(subOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i8.GSR = "ENABLED";
    FD1S3AX subOut_i9 (.D(\subOut_24__N_1135[9] ), .CK(clk_N_683), .Q(subOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i9.GSR = "ENABLED";
    FD1S3AX subOut_i10 (.D(\subOut_24__N_1135[10] ), .CK(clk_N_683), .Q(subOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i10.GSR = "ENABLED";
    FD1S3AX subOut_i11 (.D(\subOut_24__N_1135[11] ), .CK(clk_N_683), .Q(subOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i11.GSR = "ENABLED";
    FD1S3AX subOut_i12 (.D(\subOut_24__N_1135[12] ), .CK(clk_N_683), .Q(subOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i12.GSR = "ENABLED";
    FD1S3AX subOut_i13 (.D(\subOut_24__N_1135[13] ), .CK(clk_N_683), .Q(subOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i13.GSR = "ENABLED";
    FD1S3AX subOut_i14 (.D(\subOut_24__N_1135[14] ), .CK(clk_N_683), .Q(subOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i14.GSR = "ENABLED";
    FD1S3AX subOut_i15 (.D(\subOut_24__N_1135[15] ), .CK(clk_N_683), .Q(subOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i15.GSR = "ENABLED";
    FD1S3AX subOut_i16 (.D(\subOut_24__N_1135[16] ), .CK(clk_N_683), .Q(subOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i16.GSR = "ENABLED";
    FD1S3AX subOut_i17 (.D(\subOut_24__N_1135[17] ), .CK(clk_N_683), .Q(subOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i17.GSR = "ENABLED";
    FD1S3AX subOut_i18 (.D(\subOut_24__N_1135[18] ), .CK(clk_N_683), .Q(subOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i18.GSR = "ENABLED";
    FD1S3AX subOut_i19 (.D(\subOut_24__N_1135[19] ), .CK(clk_N_683), .Q(subOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i19.GSR = "ENABLED";
    FD1S3AX subOut_i20 (.D(\subOut_24__N_1135[20] ), .CK(clk_N_683), .Q(subOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i20.GSR = "ENABLED";
    FD1S3AX subOut_i21 (.D(\subOut_24__N_1135[21] ), .CK(clk_N_683), .Q(subOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i21.GSR = "ENABLED";
    FD1S3AX subOut_i23 (.D(\subOut_24__N_1135[24] ), .CK(clk_N_683), .Q(subOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam subOut_i23.GSR = "ENABLED";
    LUT4 mux_139_i12_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[11]), 
         .D(n648[11]), .Z(n678[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i11_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[10]), 
         .D(n648[10]), .Z(n678[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i28_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[27]), 
         .D(n648[27]), .Z(n678[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i15_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[14]), 
         .D(n648[14]), .Z(n678[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i16_3_lut_4_lut (.A(n21892), .B(n21867), .C(intgOut0[15]), 
         .D(n648[15]), .Z(n678[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam mux_139_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 i18374_2_lut_3_lut_4_lut_4_lut (.A(n21870), .B(n21838), .C(n21883), 
         .D(n21888), .Z(multIn2[4])) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i18374_2_lut_3_lut_4_lut_4_lut.init = 16'h1115;
    LUT4 mux_1190_i1_3_lut_4_lut (.A(n21826), .B(n42), .C(speed_set_m2[0]), 
         .D(speed_set_m3[0]), .Z(n5046)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam mux_1190_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i2_3_lut_4_lut (.A(n21826), .B(n42), .C(n21818), .D(n57), .Z(n16214)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(136[23] 137[50])
    defparam i2_3_lut_4_lut.init = 16'hfff4;
    LUT4 i13775_2_lut_rep_396_3_lut_4_lut (.A(n21834), .B(n49), .C(n42), 
         .D(n21826), .Z(n21816)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(138[23] 139[51])
    defparam i13775_2_lut_rep_396_3_lut_4_lut.init = 16'h44f4;
    LUT4 mux_1801_i4_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[3] ), 
         .D(subIn2_24__N_1301[3]), .Z(subIn2_24__N_1114[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i6_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m4[5]), .Z(n5100)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i8_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[7] ), 
         .D(subIn2_24__N_1301[7]), .Z(subIn2_24__N_1114[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i9_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[8] ), 
         .D(subIn2_24__N_1301[8]), .Z(subIn2_24__N_1114[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i17_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m4[16]), .Z(n5122)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i10_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[9] ), 
         .D(subIn2_24__N_1301[9]), .Z(subIn2_24__N_1114[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i13_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[12] ), 
         .D(subIn2_24__N_1301[12]), .Z(subIn2_24__N_1114[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13180_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[19] ), 
         .D(\speed_m2[19] ), .Z(n5)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13180_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i20_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m4[19]), .Z(n5128)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i2_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[1] ), 
         .D(\speed_m2[1] ), .Z(subIn2_24__N_1114[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i3_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[2] ), 
         .D(\speed_m2[2] ), .Z(subIn2_24__N_1114[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13600_2_lut (.A(addOut[25]), .B(n22388), .Z(backOut2_28__N_1474[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13600_2_lut.init = 16'h2222;
    LUT4 mux_1801_i5_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[4] ), 
         .D(\speed_m2[4] ), .Z(subIn2_24__N_1114[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i6_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[5] ), 
         .D(\speed_m2[5] ), .Z(subIn2_24__N_1114[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i7_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[6] ), 
         .D(\speed_m2[6] ), .Z(subIn2_24__N_1114[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13606_2_lut (.A(addOut[24]), .B(n22388), .Z(backOut3_28__N_1503[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13606_2_lut.init = 16'h2222;
    LUT4 mux_1189_i18_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m4[17]), .Z(n5124)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i11_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[10] ), 
         .D(\speed_m2[10] ), .Z(subIn2_24__N_1114[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i12_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[11] ), 
         .D(\speed_m2[11] ), .Z(subIn2_24__N_1114[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i14_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[13] ), 
         .D(\speed_m2[13] ), .Z(subIn2_24__N_1114[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13599_2_lut (.A(addOut[23]), .B(n22388), .Z(backOut2_28__N_1474[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13599_2_lut.init = 16'h2222;
    LUT4 i5_4_lut (.A(n9_c), .B(n7_adj_1836), .C(n1208[10]), .D(n1208[13]), 
         .Z(n30_adj_1819)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    CCU2D add_16120_23 (.A0(addOut[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18906), .COUT(n18907));
    defparam add_16120_23.INIT0 = 16'h0aaa;
    defparam add_16120_23.INIT1 = 16'h0aaa;
    defparam add_16120_23.INJECT1_0 = "NO";
    defparam add_16120_23.INJECT1_1 = "NO";
    LUT4 i3_2_lut (.A(n1208[14]), .B(n1208[12]), .Z(n9_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 mux_1801_i15_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[14] ), 
         .D(\speed_m2[14] ), .Z(subIn2_24__N_1114[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i16_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[15] ), 
         .D(\speed_m2[15] ), .Z(subIn2_24__N_1114[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_adj_48 (.A(n1208[11]), .B(n1208[9]), .C(n10_adj_1837), 
         .D(n1208[7]), .Z(n7_adj_1836)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_48.init = 16'haaa8;
    LUT4 mux_1801_i17_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[16] ), 
         .D(\speed_m2[16] ), .Z(subIn2_24__N_1114[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4_4_lut_adj_49 (.A(n1208[6]), .B(n8), .C(n1208[4]), .D(n4), 
         .Z(n10_adj_1837)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_49.init = 16'hfeee;
    LUT4 mux_1801_i18_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[17] ), 
         .D(\speed_m2[17] ), .Z(subIn2_24__N_1114[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1801_i19_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[18] ), 
         .D(\speed_m2[18] ), .Z(subIn2_24__N_1114[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i15_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m4[14]), .Z(n5118)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut (.A(n22388), .B(n920), .C(addOut[7]), .D(n3636), 
         .Z(intgOut1_28__N_766[7])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1110;
    LUT4 i2_2_lut_adj_50 (.A(n1208[5]), .B(n1208[8]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_50.init = 16'heeee;
    LUT4 i1_4_lut_adj_51 (.A(n1208[3]), .B(n1208[2]), .C(n1208[1]), .D(n1208[0]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_51.init = 16'haaa8;
    LUT4 mux_1801_i1_3_lut_4_lut (.A(ss[2]), .B(n21877), .C(\speed_m1[0] ), 
         .D(\speed_m2[0] ), .Z(subIn2_24__N_1114[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1801_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i5_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m4[4]), .Z(n5098)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut_adj_52 (.A(n22388), .B(n920), .C(addOut[8]), .D(n3636), 
         .Z(intgOut0_28__N_735[8])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_52.init = 16'h1110;
    PFUMX i18450 (.BLUT(n21925), .ALUT(n21926), .C0(n22388), .Z(clk_N_683_enable_240));
    LUT4 mux_138_i22_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[21]), 
         .D(intgOut2[21]), .Z(n648[21])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i22_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i28_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[27]), 
         .D(intgOut2[27]), .Z(n648[27])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i28_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i20_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[19]), 
         .D(intgOut2[19]), .Z(n648[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i20_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i11_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[10]), 
         .D(intgOut2[10]), .Z(n648[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i29_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[28]), 
         .D(intgOut2[28]), .Z(n648[28])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i29_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i9_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[8]), 
         .D(intgOut2[8]), .Z(n648[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i9_3_lut_4_lut.init = 16'hfe10;
    LUT4 i53_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[0]), .D(intgOut2[0]), 
         .Z(n28)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam i53_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13598_2_lut (.A(addOut[22]), .B(n22388), .Z(backOut2_28__N_1474[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13598_2_lut.init = 16'h2222;
    LUT4 mux_138_i14_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[13]), 
         .D(intgOut2[13]), .Z(n648[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i14_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_4_lut_adj_53 (.A(n22388), .B(n920), .C(addOut[10]), 
         .D(n3636), .Z(intgOut0_28__N_735[10])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_53.init = 16'h1110;
    LUT4 mux_1189_i10_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m4[9]), .Z(n5108)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i25_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[24]), 
         .D(intgOut2[24]), .Z(n648[24])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 i41_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[3]), .D(intgOut2[3]), 
         .Z(n23)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam i41_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i8_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[7]), 
         .D(intgOut2[7]), .Z(n648[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i18_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[17]), 
         .D(intgOut2[17]), .Z(n648[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i18_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1189_i13_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m4[12]), .Z(n5114)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i13_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_16120_21 (.A0(addOut[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18905), .COUT(n18906));
    defparam add_16120_21.INIT0 = 16'h0aaa;
    defparam add_16120_21.INIT1 = 16'h0aaa;
    defparam add_16120_21.INJECT1_0 = "NO";
    defparam add_16120_21.INJECT1_1 = "NO";
    CCU2D add_16120_19 (.A0(addOut[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18904), .COUT(n18905));
    defparam add_16120_19.INIT0 = 16'hf555;
    defparam add_16120_19.INIT1 = 16'hf555;
    defparam add_16120_19.INJECT1_0 = "NO";
    defparam add_16120_19.INJECT1_1 = "NO";
    LUT4 i5_4_lut_adj_54 (.A(n9_adj_1838), .B(n7_adj_1839), .C(n1187[10]), 
         .D(n1187[13]), .Z(n30_adj_1818)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_54.init = 16'h8000;
    LUT4 i3_2_lut_adj_55 (.A(n1187[14]), .B(n1187[12]), .Z(n9_adj_1838)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_55.init = 16'h8888;
    LUT4 i1_4_lut_adj_56 (.A(n1187[11]), .B(n1187[9]), .C(n10_adj_1840), 
         .D(n1187[7]), .Z(n7_adj_1839)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_56.init = 16'haaa8;
    LUT4 i4_4_lut_adj_57 (.A(n1187[6]), .B(n8_adj_1841), .C(n1187[4]), 
         .D(n4_adj_1842), .Z(n10_adj_1840)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_57.init = 16'hfeee;
    LUT4 i2_2_lut_adj_58 (.A(n1187[5]), .B(n1187[8]), .Z(n8_adj_1841)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_58.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_59 (.A(n22388), .B(n920), .C(addOut[11]), 
         .D(n3636), .Z(intgOut1_28__N_766[11])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_59.init = 16'h1110;
    LUT4 i1_4_lut_adj_60 (.A(n1187[3]), .B(n1187[2]), .C(n1187[1]), .D(n1187[0]), 
         .Z(n4_adj_1842)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_60.init = 16'haaa8;
    LUT4 mux_138_i26_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[25]), 
         .D(intgOut2[25]), .Z(n648[25])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i26_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i7_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[6]), 
         .D(intgOut2[6]), .Z(n648[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 i41_3_lut_4_lut_adj_61 (.A(n21888), .B(n21869), .C(intgOut1[2]), 
         .D(intgOut2[2]), .Z(n23_adj_1829)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam i41_3_lut_4_lut_adj_61.init = 16'hfe10;
    LUT4 i1_3_lut_4_lut_adj_62 (.A(n22388), .B(n920), .C(addOut[12]), 
         .D(n3636), .Z(intgOut1_28__N_766[12])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_62.init = 16'h1110;
    LUT4 mux_1189_i11_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m4[10]), .Z(n5110)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i41_3_lut_4_lut_adj_63 (.A(n21888), .B(n21869), .C(intgOut1[5]), 
         .D(intgOut2[5]), .Z(n23_adj_1833)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam i41_3_lut_4_lut_adj_63.init = 16'hfe10;
    LUT4 mux_138_i10_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[9]), 
         .D(intgOut2[9]), .Z(n648[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i10_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1189_i9_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m4[8]), .Z(n5106)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i21_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[20]), 
         .D(intgOut2[20]), .Z(n648[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i23_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[22]), 
         .D(intgOut2[22]), .Z(n648[22])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i23_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_179_17 (.A0(Out0[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18689), 
          .S0(n1145[15]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_17.INIT0 = 16'h5aaa;
    defparam add_179_17.INIT1 = 16'h0000;
    defparam add_179_17.INJECT1_0 = "NO";
    defparam add_179_17.INJECT1_1 = "NO";
    LUT4 mux_1189_i8_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m4[7]), .Z(n5104)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i7_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m4[6]), .Z(n5102)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i24_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[23]), 
         .D(intgOut2[23]), .Z(n648[23])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i24_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_16120_17 (.A0(addOut[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18903), .COUT(n18904));
    defparam add_16120_17.INIT0 = 16'hf555;
    defparam add_16120_17.INIT1 = 16'hf555;
    defparam add_16120_17.INJECT1_0 = "NO";
    defparam add_16120_17.INJECT1_1 = "NO";
    LUT4 mux_1189_i1_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m4[0]), .Z(n5048)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i27_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[26]), 
         .D(intgOut2[26]), .Z(n648[26])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i27_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i17_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[16]), 
         .D(intgOut2[16]), .Z(n648[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i17_3_lut_4_lut.init = 16'hfe10;
    LUT4 i41_3_lut_4_lut_adj_64 (.A(n21888), .B(n21869), .C(intgOut1[1]), 
         .D(intgOut2[1]), .Z(n23_adj_1831)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam i41_3_lut_4_lut_adj_64.init = 16'hfe10;
    LUT4 mux_1189_i2_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m4[1]), .Z(n5092)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i19_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[18]), 
         .D(intgOut2[18]), .Z(n648[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i19_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i13_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[12]), 
         .D(intgOut2[12]), .Z(n648[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 i41_3_lut_4_lut_adj_65 (.A(n21888), .B(n21869), .C(intgOut1[4]), 
         .D(intgOut2[4]), .Z(n23_adj_1827)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam i41_3_lut_4_lut_adj_65.init = 16'hfe10;
    LUT4 mux_138_i12_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[11]), 
         .D(intgOut2[11]), .Z(n648[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i12_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i15_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[14]), 
         .D(intgOut2[14]), .Z(n648[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i16_3_lut_4_lut (.A(n21888), .B(n21869), .C(intgOut1[15]), 
         .D(intgOut2[15]), .Z(n648[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(169[9:16])
    defparam mux_138_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1189_i19_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m4[18]), .Z(n5126)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i19_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX dutyout_m4_i0_i9 (.D(n1390[9]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i8 (.D(n1390[8]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i7 (.D(n1390[7]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i6 (.D(n1390[6]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i5 (.D(n1390[5]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i4 (.D(n2189[4]), .SP(clk_N_683_enable_392), .CD(n13107), 
            .CK(clk_N_683), .Q(PWMdut_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i3 (.D(n1390[3]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i2 (.D(n2189[2]), .SP(clk_N_683_enable_392), .CD(n13107), 
            .CK(clk_N_683), .Q(PWMdut_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i1 (.D(n2189[1]), .SP(clk_N_683_enable_392), .CD(n13107), 
            .CK(clk_N_683), .Q(PWMdut_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i9 (.D(n1346[9]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i8 (.D(n1346[8]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i7 (.D(n1346[7]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i6 (.D(n1346[6]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i5 (.D(n1346[5]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i5.GSR = "DISABLED";
    CCU2D add_179_15 (.A0(Out0[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18688), 
          .COUT(n18689), .S0(n1145[13]), .S1(n1145[14]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_15.INIT0 = 16'h5aaa;
    defparam add_179_15.INIT1 = 16'h5aaa;
    defparam add_179_15.INJECT1_0 = "NO";
    defparam add_179_15.INJECT1_1 = "NO";
    LUT4 mux_1189_i14_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m4[13]), .Z(n5116)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i4_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m4[3]), .Z(n5096)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i4_3_lut (.A(\speed_m3[3] ), .B(\speed_m2[3] ), .C(n22376), 
         .Z(subIn2_24__N_1301[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i4_3_lut.init = 16'hcaca;
    LUT4 i18315_3_lut_3_lut_4_lut_4_lut (.A(n21892), .B(n21869), .C(n21858), 
         .D(n21867), .Z(n20525)) /* synthesis lut_function=(!(A (B (C (D)))+!A (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(170[9:16])
    defparam i18315_3_lut_3_lut_4_lut_4_lut.init = 16'h2faf;
    LUT4 i1_2_lut_3_lut_4_lut_adj_66 (.A(n920), .B(n3636), .C(addOut[5]), 
         .D(n22388), .Z(intgOut1_28__N_766[5])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_66.init = 16'h0010;
    LUT4 mux_1189_i3_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m4[2]), .Z(n5094)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i16_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m4[15]), .Z(n5120)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i21_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m4[20]), .Z(n5130)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_4_lut (.A(n21885), .B(n22388), .C(n20247), .D(n21903), 
         .Z(clk_N_683_enable_268)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B+((D)+!C))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h88b8;
    LUT4 mux_1189_i12_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m4[11]), .Z(n5112)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(134[23] 135[50])
    defparam mux_1189_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_4_lut_adj_67 (.A(n21885), .B(n22388), .C(n20202), .D(ss[1]), 
         .Z(clk_N_683_enable_184)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(B+(C+!(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_67.init = 16'h8b88;
    LUT4 i1_4_lut_4_lut_adj_68 (.A(n21885), .B(n22388), .C(n20199), .D(n21903), 
         .Z(clk_N_683_enable_212)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+(C+(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_68.init = 16'h888b;
    LUT4 i1_4_lut_4_lut_adj_69 (.A(n21885), .B(n22388), .C(n20202), .D(ss[1]), 
         .Z(clk_N_683_enable_156)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+(C+(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_69.init = 16'h888b;
    LUT4 mux_1800_i8_3_lut (.A(\speed_m3[7] ), .B(\speed_m2[7] ), .C(n22376), 
         .Z(subIn2_24__N_1301[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_70 (.A(n21885), .B(n22388), .C(n21884), .D(ss[3]), 
         .Z(clk_N_683_enable_296)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_70.init = 16'hb888;
    LUT4 mux_1800_i9_3_lut (.A(\speed_m3[8] ), .B(\speed_m2[8] ), .C(n22376), 
         .Z(subIn2_24__N_1301[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i9_3_lut.init = 16'hcaca;
    LUT4 i13597_2_lut (.A(addOut[21]), .B(n22388), .Z(backOut2_28__N_1474[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13597_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_adj_71 (.A(n22388), .B(n920), .C(addOut[13]), 
         .D(n3636), .Z(intgOut1_28__N_766[13])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_71.init = 16'h1110;
    LUT4 mux_1800_i10_3_lut (.A(\speed_m3[9] ), .B(\speed_m2[9] ), .C(n22376), 
         .Z(subIn2_24__N_1301[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i10_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_72 (.A(n22388), .B(n920), .C(addOut[15]), 
         .D(n3636), .Z(intgOut2_28__N_795[15])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_72.init = 16'h1110;
    LUT4 mux_1800_i13_3_lut (.A(\speed_m3[12] ), .B(\speed_m2[12] ), .C(n22376), 
         .Z(subIn2_24__N_1301[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1800_i2_4_lut (.A(\speed_m4[1] ), .B(\speed_m3[1] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i2_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i3_4_lut (.A(\speed_m4[2] ), .B(\speed_m3[2] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i3_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i5_4_lut (.A(\speed_m4[4] ), .B(\speed_m3[4] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i5_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_4_lut_adj_73 (.A(n22388), .B(n920), .C(addOut[20]), 
         .D(n3636), .Z(intgOut1_28__N_766[20])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_73.init = 16'h1110;
    LUT4 mux_1800_i6_4_lut (.A(\speed_m4[5] ), .B(\speed_m3[5] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i6_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_4_lut_adj_74 (.A(n22388), .B(n920), .C(addOut[21]), 
         .D(n3636), .Z(intgOut1_28__N_766[21])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_74.init = 16'h1110;
    LUT4 mux_1800_i7_4_lut (.A(\speed_m4[6] ), .B(\speed_m3[6] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i7_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i11_4_lut (.A(\speed_m4[10] ), .B(\speed_m3[10] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i11_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i12_4_lut (.A(\speed_m4[11] ), .B(\speed_m3[11] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i12_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i14_4_lut (.A(\speed_m4[13] ), .B(\speed_m3[13] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i14_4_lut.init = 16'hcac0;
    LUT4 i13566_4_lut_4_lut (.A(n920), .B(n3636), .C(addOut[9]), .D(n22388), 
         .Z(intgOut1_28__N_766[9])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13566_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_1800_i15_4_lut (.A(\speed_m4[14] ), .B(\speed_m3[14] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i15_4_lut.init = 16'hcac0;
    LUT4 i5_4_lut_adj_75 (.A(n9_adj_1843), .B(n7_adj_1844), .C(n1166[10]), 
         .D(n1166[13]), .Z(n30_c)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_75.init = 16'h8000;
    LUT4 mux_1800_i16_4_lut (.A(\speed_m4[15] ), .B(\speed_m3[15] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i16_4_lut.init = 16'hcac0;
    LUT4 i3_2_lut_adj_76 (.A(n1166[14]), .B(n1166[12]), .Z(n9_adj_1843)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_76.init = 16'h8888;
    LUT4 i1_4_lut_adj_77 (.A(n1166[11]), .B(n1166[9]), .C(n10_adj_1845), 
         .D(n1166[7]), .Z(n7_adj_1844)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_77.init = 16'haaa8;
    LUT4 i4_4_lut_adj_78 (.A(n1166[6]), .B(n8_adj_1846), .C(n1166[4]), 
         .D(n4_adj_1847), .Z(n10_adj_1845)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_78.init = 16'hfeee;
    LUT4 i2_2_lut_adj_79 (.A(n1166[5]), .B(n1166[8]), .Z(n8_adj_1846)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_79.init = 16'heeee;
    LUT4 i1_4_lut_adj_80 (.A(n1166[3]), .B(n1166[2]), .C(n1166[1]), .D(n1166[0]), 
         .Z(n4_adj_1847)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_80.init = 16'haaa8;
    LUT4 mux_1800_i17_4_lut (.A(\speed_m4[16] ), .B(\speed_m3[16] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i17_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i18_4_lut (.A(\speed_m4[17] ), .B(\speed_m3[17] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i18_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i19_4_lut (.A(\speed_m4[18] ), .B(\speed_m3[18] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i19_4_lut.init = 16'hcac0;
    LUT4 mux_1800_i1_4_lut (.A(\speed_m4[0] ), .B(\speed_m3[0] ), .C(n21857), 
         .D(n4133), .Z(subIn2_24__N_1301[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(147[18] 151[17])
    defparam mux_1800_i1_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_4_lut_adj_81 (.A(n22388), .B(n920), .C(addOut[22]), 
         .D(n3636), .Z(intgOut2_28__N_795[22])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_81.init = 16'h1110;
    LUT4 mux_1245_i2_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[1]), 
         .D(speed_set_m4[1]), .Z(n2485[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i2_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i13_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[12]), 
         .D(speed_set_m4[12]), .Z(n2485[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i16_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[15]), 
         .D(speed_set_m4[15]), .Z(n2485[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i17_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[16]), 
         .D(speed_set_m4[16]), .Z(n2485[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i17_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_4_lut_adj_82 (.A(n22388), .B(n920), .C(addOut[23]), 
         .D(n3636), .Z(intgOut1_28__N_766[23])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_82.init = 16'h1110;
    CCU2D add_16120_15 (.A0(addOut[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18902), .COUT(n18903));
    defparam add_16120_15.INIT0 = 16'hf555;
    defparam add_16120_15.INIT1 = 16'h0aaa;
    defparam add_16120_15.INJECT1_0 = "NO";
    defparam add_16120_15.INJECT1_1 = "NO";
    CCU2D add_16120_13 (.A0(addOut[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18901), .COUT(n18902));
    defparam add_16120_13.INIT0 = 16'h0aaa;
    defparam add_16120_13.INIT1 = 16'h0aaa;
    defparam add_16120_13.INJECT1_0 = "NO";
    defparam add_16120_13.INJECT1_1 = "NO";
    LUT4 mux_1245_i18_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[17]), 
         .D(speed_set_m4[17]), .Z(n2485[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i18_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i5_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[4]), 
         .D(speed_set_m4[4]), .Z(n2485[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i5_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_16120_11 (.A0(addOut[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18900), .COUT(n18901));
    defparam add_16120_11.INIT0 = 16'h0aaa;
    defparam add_16120_11.INIT1 = 16'h0aaa;
    defparam add_16120_11.INJECT1_0 = "NO";
    defparam add_16120_11.INJECT1_1 = "NO";
    LUT4 i13587_2_lut (.A(addOut[20]), .B(n22388), .Z(backOut1_28__N_1445[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13587_2_lut.init = 16'h2222;
    LUT4 mux_1245_i3_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[2]), 
         .D(speed_set_m4[2]), .Z(n2485[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i11_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[10]), 
         .D(speed_set_m4[10]), .Z(n2485[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 ss_1__bdd_4_lut (.A(n22388), .B(ss[0]), .C(ss[2]), .D(ss[3]), 
         .Z(n16286)) /* synthesis lut_function=(A+(B+(C (D)+!C !(D)))) */ ;
    defparam ss_1__bdd_4_lut.init = 16'hfeef;
    LUT4 mux_1245_i6_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[5]), 
         .D(speed_set_m4[5]), .Z(n2485[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_4_lut_adj_83 (.A(n22388), .B(n920), .C(addOut[24]), 
         .D(n3636), .Z(intgOut0_28__N_735[24])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_83.init = 16'h1110;
    LUT4 i1_3_lut_4_lut_adj_84 (.A(n22388), .B(n920), .C(addOut[25]), 
         .D(n3636), .Z(intgOut1_28__N_766[25])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_84.init = 16'h1110;
    LUT4 mux_1245_i7_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[6]), 
         .D(speed_set_m4[6]), .Z(n2485[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i7_3_lut_4_lut.init = 16'hfe10;
    FD1P3IX dutyout_m3_i0_i4 (.D(n2177[4]), .SP(clk_N_683_enable_392), .CD(n13098), 
            .CK(clk_N_683), .Q(PWMdut_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i3 (.D(n1346[3]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i2 (.D(n2177[2]), .SP(clk_N_683_enable_392), .CD(n13098), 
            .CK(clk_N_683), .Q(PWMdut_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i1 (.D(n2177[1]), .SP(clk_N_683_enable_392), .CD(n13098), 
            .CK(clk_N_683), .Q(PWMdut_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i9 (.D(n1302[9]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i8 (.D(n1302[8]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i8.GSR = "DISABLED";
    LUT4 mux_135_i25_4_lut (.A(backOut2_c[24]), .B(backOut3_c[24]), .C(n21851), 
         .D(n9), .Z(n558[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i25_4_lut.init = 16'h0aca;
    LUT4 mux_1245_i19_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[18]), 
         .D(speed_set_m4[18]), .Z(n2485[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i19_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i17_4_lut (.A(backOut2_c[16]), .B(backOut3_c[16]), .C(n21851), 
         .D(n9), .Z(n558[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i17_4_lut.init = 16'h0aca;
    LUT4 i13586_2_lut (.A(addOut[19]), .B(n22388), .Z(backOut1_28__N_1445[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13586_2_lut.init = 16'h2222;
    LUT4 i13755_2_lut (.A(addOut[18]), .B(n22388), .Z(backOut2_28__N_1474[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13755_2_lut.init = 16'h2222;
    CCU2D add_16120_9 (.A0(addOut[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18899), .COUT(n18900));
    defparam add_16120_9.INIT0 = 16'h0aaa;
    defparam add_16120_9.INIT1 = 16'hf555;
    defparam add_16120_9.INJECT1_0 = "NO";
    defparam add_16120_9.INJECT1_1 = "NO";
    LUT4 mux_1245_i15_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[14]), 
         .D(speed_set_m4[14]), .Z(n2485[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i4_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[3]), 
         .D(speed_set_m4[3]), .Z(n2485[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i1_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[0]), 
         .D(speed_set_m4[0]), .Z(n2485[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i7_4_lut (.A(backOut2_c[6]), .B(backOut3_c[6]), .C(n21851), 
         .D(n9), .Z(n558[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i7_4_lut.init = 16'h0aca;
    LUT4 mux_1245_i21_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[20]), 
         .D(speed_set_m4[20]), .Z(n2485[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i21_3_lut_4_lut.init = 16'hfe10;
    FD1P3IX dutyout_m2_i0_i7 (.D(n1302[7]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i6 (.D(n1302[6]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i5 (.D(n1302[5]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i4 (.D(n2165[4]), .SP(clk_N_683_enable_392), .CD(n13089), 
            .CK(clk_N_683), .Q(PWMdut_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i3 (.D(n1302[3]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i2 (.D(n2165[2]), .SP(clk_N_683_enable_392), .CD(n13089), 
            .CK(clk_N_683), .Q(PWMdut_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i2.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_85 (.A(n22388), .B(n920), .C(addOut[26]), 
         .D(n3636), .Z(intgOut1_28__N_766[26])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_85.init = 16'h1110;
    LUT4 mux_1245_i8_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[7]), 
         .D(speed_set_m4[7]), .Z(n2485[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i26_4_lut (.A(backOut2_c[25]), .B(backOut3_c[25]), .C(n21851), 
         .D(n9), .Z(n558[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i26_4_lut.init = 16'h0aca;
    LUT4 mux_1245_i20_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[19]), 
         .D(speed_set_m4[19]), .Z(n2485[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i20_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i18_4_lut (.A(backOut2_c[17]), .B(backOut3_c[17]), .C(n21851), 
         .D(n9), .Z(n558[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i18_4_lut.init = 16'h0aca;
    FD1P3IX dutyout_m4_i0_i0 (.D(n2189[0]), .SP(clk_N_683_enable_392), .CD(n13107), 
            .CK(clk_N_683), .Q(PWMdut_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i0.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i0 (.D(n2177[0]), .SP(clk_N_683_enable_392), .CD(n13098), 
            .CK(clk_N_683), .Q(PWMdut_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i0.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i0 (.D(n2165[0]), .SP(clk_N_683_enable_392), .CD(n13089), 
            .CK(clk_N_683), .Q(PWMdut_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i0.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i0 (.D(n2153[0]), .SP(clk_N_683_enable_392), .CD(n13080), 
            .CK(clk_N_683), .Q(PWMdut_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i0.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i1 (.D(n2165[1]), .SP(clk_N_683_enable_392), .CD(n13089), 
            .CK(clk_N_683), .Q(PWMdut_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i9 (.D(n1258[9]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i8 (.D(n1258[8]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i7 (.D(n1258[7]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i6 (.D(n1258[6]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i5 (.D(n1258[5]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i5.GSR = "DISABLED";
    LUT4 i13750_2_lut (.A(addOut[17]), .B(n22388), .Z(backOut3_28__N_1503[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13750_2_lut.init = 16'h2222;
    FD1P3IX dutyout_m1_i0_i4 (.D(n2153[4]), .SP(clk_N_683_enable_392), .CD(n13080), 
            .CK(clk_N_683), .Q(PWMdut_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i3 (.D(n1258[3]), .SP(clk_N_683_enable_392), .CD(n13082), 
            .CK(clk_N_683), .Q(PWMdut_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i2 (.D(n2153[2]), .SP(clk_N_683_enable_392), .CD(n13080), 
            .CK(clk_N_683), .Q(PWMdut_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i1 (.D(n2153[1]), .SP(clk_N_683_enable_392), .CD(n13080), 
            .CK(clk_N_683), .Q(PWMdut_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i1.GSR = "DISABLED";
    LUT4 mux_1245_i9_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[8]), 
         .D(speed_set_m4[8]), .Z(n2485[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i9_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i8_4_lut (.A(backOut2_c[7]), .B(backOut3_c[7]), .C(n21851), 
         .D(n9), .Z(n558[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i8_4_lut.init = 16'h0aca;
    LUT4 mux_1245_i10_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[9]), 
         .D(speed_set_m4[9]), .Z(n2485[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i10_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_4_lut_adj_86 (.A(n22388), .B(n920), .C(addOut[27]), 
         .D(n3636), .Z(intgOut1_28__N_766[27])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_86.init = 16'h1110;
    LUT4 i1_2_lut_adj_87 (.A(ss[1]), .B(ss[2]), .Z(n20199)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_adj_87.init = 16'hbbbb;
    LUT4 mux_1245_i14_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[13]), 
         .D(speed_set_m4[13]), .Z(n2485[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i14_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1245_i12_3_lut_4_lut (.A(n21834), .B(n49), .C(speed_set_m3[11]), 
         .D(speed_set_m4[11]), .Z(n2485[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1245_i12_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3410_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m2[10]), .Z(n5707)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3410_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_179_13 (.A0(Out0[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18687), 
          .COUT(n18688), .S0(n1145[11]), .S1(n1145[12]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_13.INIT0 = 16'h5aaa;
    defparam add_179_13.INIT1 = 16'h5aaa;
    defparam add_179_13.INJECT1_0 = "NO";
    defparam add_179_13.INJECT1_1 = "NO";
    LUT4 i18319_2_lut_rep_395_2_lut_3_lut_4_lut (.A(n21824), .B(n35), .C(n42), 
         .D(n21826), .Z(n21815)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))))) */ ;
    defparam i18319_2_lut_rep_395_2_lut_3_lut_4_lut.init = 16'h111f;
    LUT4 i3392_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m2[1]), .Z(n5689)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3392_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3394_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m2[2]), .Z(n5691)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3394_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i27_4_lut (.A(backOut2_c[26]), .B(backOut3_c[26]), .C(n21851), 
         .D(n9), .Z(n558[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i27_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_88 (.A(n920), .B(n3636), .C(addOut[0]), 
         .D(n22388), .Z(intgOut0_28__N_735[0])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_88.init = 16'h0010;
    LUT4 i1_3_lut_4_lut_adj_89 (.A(n22388), .B(n920), .C(addOut[28]), 
         .D(n3636), .Z(intgOut1_28__N_766[28])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_89.init = 16'h1110;
    LUT4 i3396_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m2[3]), .Z(n5693)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3396_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3398_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m2[4]), .Z(n5695)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3398_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3400_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m2[5]), .Z(n5697)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3400_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i19_4_lut (.A(backOut2_c[18]), .B(backOut3_c[18]), .C(n21851), 
         .D(n9), .Z(n558[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i19_4_lut.init = 16'h0aca;
    LUT4 i13756_2_lut (.A(addOut[16]), .B(n22388), .Z(backOut2_28__N_1474[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13756_2_lut.init = 16'h2222;
    CCU2D add_16120_7 (.A0(addOut[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18898), .COUT(n18899));
    defparam add_16120_7.INIT0 = 16'h0aaa;
    defparam add_16120_7.INIT1 = 16'h0aaa;
    defparam add_16120_7.INJECT1_0 = "NO";
    defparam add_16120_7.INJECT1_1 = "NO";
    CCU2D add_179_11 (.A0(Out0[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18686), 
          .COUT(n18687), .S0(n1145[9]), .S1(n1145[10]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_11.INIT0 = 16'h5aaa;
    defparam add_179_11.INIT1 = 16'h5aaa;
    defparam add_179_11.INJECT1_0 = "NO";
    defparam add_179_11.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_90 (.A(n21818), .B(n21817), .C(n21839), .D(n21819), 
         .Z(n7_c)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i2_3_lut_4_lut_adj_90.init = 16'hffef;
    LUT4 i17423_2_lut (.A(ss[2]), .B(ss[1]), .Z(n20247)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17423_2_lut.init = 16'h8888;
    LUT4 i3402_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m2[6]), .Z(n5699)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3402_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i9_4_lut (.A(backOut2_c[8]), .B(backOut3_c[8]), .C(n21851), 
         .D(n9), .Z(n558[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i9_4_lut.init = 16'h0aca;
    LUT4 i13757_2_lut (.A(addOut[15]), .B(n22388), .Z(backOut2_28__N_1474[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13757_2_lut.init = 16'h2222;
    LUT4 i3404_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m2[7]), .Z(n5701)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3404_3_lut_4_lut.init = 16'hfe10;
    LUT4 i5_4_lut_adj_91 (.A(n9_adj_1849), .B(n7_adj_1850), .C(n1145[10]), 
         .D(n1145[13]), .Z(n30_adj_1851)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_91.init = 16'h8000;
    LUT4 i3_2_lut_adj_92 (.A(n1145[14]), .B(n1145[12]), .Z(n9_adj_1849)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_92.init = 16'h8888;
    LUT4 mux_135_i28_4_lut (.A(backOut2_c[27]), .B(backOut3_c[27]), .C(n21851), 
         .D(n9), .Z(n558[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i28_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_93 (.A(n1145[11]), .B(n1145[9]), .C(n10_adj_1852), 
         .D(n1145[7]), .Z(n7_adj_1850)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_93.init = 16'haaa8;
    CCU2D add_16120_5 (.A0(addOut[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18897), .COUT(n18898));
    defparam add_16120_5.INIT0 = 16'hf555;
    defparam add_16120_5.INIT1 = 16'hf555;
    defparam add_16120_5.INJECT1_0 = "NO";
    defparam add_16120_5.INJECT1_1 = "NO";
    LUT4 i4_4_lut_adj_94 (.A(n1145[6]), .B(n8_adj_1853), .C(n1145[4]), 
         .D(n4_adj_1854), .Z(n10_adj_1852)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_94.init = 16'hfeee;
    LUT4 i2_2_lut_adj_95 (.A(n1145[5]), .B(n1145[8]), .Z(n8_adj_1853)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_95.init = 16'heeee;
    LUT4 i1_4_lut_adj_96 (.A(n1145[3]), .B(n1145[2]), .C(n1145[1]), .D(n1145[0]), 
         .Z(n4_adj_1854)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_96.init = 16'haaa8;
    LUT4 i3406_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m2[8]), .Z(n5703)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3406_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i20_4_lut (.A(backOut2_c[19]), .B(backOut3_c[19]), .C(n21851), 
         .D(n9), .Z(n558[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i20_4_lut.init = 16'h0aca;
    CCU2D add_16120_3 (.A0(addOut[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18896), .COUT(n18897));
    defparam add_16120_3.INIT0 = 16'hf555;
    defparam add_16120_3.INIT1 = 16'hf555;
    defparam add_16120_3.INJECT1_0 = "NO";
    defparam add_16120_3.INJECT1_1 = "NO";
    LUT4 i7_4_lut_adj_97 (.A(Out3[3]), .B(n14_adj_1855), .C(n10_adj_1856), 
         .D(Out3[4]), .Z(n19124)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam i7_4_lut_adj_97.init = 16'hfffe;
    LUT4 i6_4_lut_adj_98 (.A(Out3[11]), .B(Out3[7]), .C(Out3[2]), .D(Out3[10]), 
         .Z(n14_adj_1855)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam i6_4_lut_adj_98.init = 16'hfffe;
    LUT4 i2_2_lut_adj_99 (.A(Out3[9]), .B(Out3[1]), .Z(n10_adj_1856)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam i2_2_lut_adj_99.init = 16'heeee;
    LUT4 i4_4_lut_adj_100 (.A(Out3[5]), .B(Out3[6]), .C(Out3[0]), .D(n6_adj_1857), 
         .Z(n19125)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam i4_4_lut_adj_100.init = 16'hfffe;
    LUT4 i1_2_lut_adj_101 (.A(Out3[8]), .B(Out3[12]), .Z(n6_adj_1857)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam i1_2_lut_adj_101.init = 16'heeee;
    LUT4 i1_2_lut_4_lut (.A(n22388), .B(n21922), .C(ss[3]), .D(ss[0]), 
         .Z(multIn2[6])) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h1400;
    LUT4 i2_3_lut_4_lut_adj_102 (.A(ss[2]), .B(n21898), .C(n22388), .D(ss[1]), 
         .Z(n20197)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i2_3_lut_4_lut_adj_102.init = 16'h0800;
    CCU2D add_16120_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[0]), .B1(addOut[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18896));
    defparam add_16120_1.INIT0 = 16'hF000;
    defparam add_16120_1.INIT1 = 16'ha666;
    defparam add_16120_1.INJECT1_0 = "NO";
    defparam add_16120_1.INJECT1_1 = "NO";
    LUT4 i18261_2_lut_3_lut_4_lut (.A(n21893), .B(n22375), .C(n22376), 
         .D(ss[2]), .Z(n20586)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i18261_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i13758_2_lut (.A(addOut[14]), .B(n22388), .Z(backOut2_28__N_1474[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13758_2_lut.init = 16'h2222;
    LUT4 i3408_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m2[9]), .Z(n5705)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3408_3_lut_4_lut.init = 16'hfe10;
    LUT4 n11061_bdd_4_lut_rep_506 (.A(n21893), .B(ss[0]), .C(n22379), 
         .D(ss[1]), .Z(n22376)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam n11061_bdd_4_lut_rep_506.init = 16'h0410;
    LUT4 i13585_2_lut (.A(addOut[13]), .B(n22388), .Z(backOut1_28__N_1445[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13585_2_lut.init = 16'h2222;
    LUT4 i3412_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m2[11]), .Z(n5709)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3412_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3414_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m2[12]), .Z(n5711)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3414_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_179_9 (.A0(Out0[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18685), 
          .COUT(n18686), .S0(n1145[7]), .S1(n1145[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_9.INIT0 = 16'h5aaa;
    defparam add_179_9.INIT1 = 16'h5aaa;
    defparam add_179_9.INJECT1_0 = "NO";
    defparam add_179_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_103 (.A(n21923), .B(n21922), .C(n22383), 
         .D(n22388), .Z(n20184)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_3_lut_4_lut_adj_103.init = 16'he0f0;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n21923), .B(n21922), .C(n20247), .D(n22388), 
         .Z(clk_N_683_enable_128)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_4_lut_4_lut_4_lut.init = 16'hee50;
    LUT4 i1_4_lut_4_lut_4_lut_adj_104 (.A(n21923), .B(n21922), .C(n20199), 
         .D(n22388), .Z(clk_N_683_enable_100)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_4_lut_4_lut_4_lut_adj_104.init = 16'hee05;
    LUT4 i13769_2_lut_rep_466 (.A(ss[1]), .B(ss[3]), .Z(n21886)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13769_2_lut_rep_466.init = 16'heeee;
    LUT4 i2_3_lut_4_lut_adj_105 (.A(ss[1]), .B(ss[3]), .C(n22379), .D(ss[0]), 
         .Z(n19129)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_105.init = 16'hfffe;
    LUT4 i3416_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m2[13]), .Z(n5713)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3416_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3418_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m2[14]), .Z(n5715)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3418_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_179_7 (.A0(Out0[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18684), 
          .COUT(n18685), .S0(n1145[5]), .S1(n1145[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_7.INIT0 = 16'h5aaa;
    defparam add_179_7.INIT1 = 16'h5aaa;
    defparam add_179_7.INJECT1_0 = "NO";
    defparam add_179_7.INJECT1_1 = "NO";
    LUT4 mux_135_i10_4_lut (.A(backOut2_c[9]), .B(backOut3_c[9]), .C(n21851), 
         .D(n9), .Z(n558[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i10_4_lut.init = 16'h0aca;
    LUT4 equal_114_i6_2_lut_rep_468 (.A(ss[0]), .B(ss[1]), .Z(n21888)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(175[9:17])
    defparam equal_114_i6_2_lut_rep_468.init = 16'hdddd;
    CCU2D add_179_5 (.A0(Out0[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18683), 
          .COUT(n18684), .S0(n1145[3]), .S1(n1145[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_5.INIT0 = 16'h5aaa;
    defparam add_179_5.INIT1 = 16'h5aaa;
    defparam add_179_5.INJECT1_0 = "NO";
    defparam add_179_5.INJECT1_1 = "NO";
    LUT4 i3420_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m2[15]), .Z(n5717)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3420_3_lut_4_lut.init = 16'hfe10;
    LUT4 i18406_2_lut_rep_415_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21894), 
         .D(n22379), .Z(n21835)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(175[9:17])
    defparam i18406_2_lut_rep_415_2_lut_3_lut_4_lut.init = 16'h0002;
    CCU2D add_179_3 (.A0(Out0[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18682), 
          .COUT(n18683), .S0(n1145[1]), .S1(n1145[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_3.INIT0 = 16'h5aaa;
    defparam add_179_3.INIT1 = 16'h5aaa;
    defparam add_179_3.INJECT1_0 = "NO";
    defparam add_179_3.INJECT1_1 = "NO";
    LUT4 i3422_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m2[16]), .Z(n5719)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3422_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3424_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m2[17]), .Z(n5721)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3424_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i11_4_lut (.A(backOut2_c[10]), .B(backOut3_c[10]), .C(n21851), 
         .D(n9), .Z(n558[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i11_4_lut.init = 16'h0aca;
    LUT4 ss_4__I_0_319_i9_2_lut_rep_438_3_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21893), .D(ss[2]), .Z(n21858)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(175[9:17])
    defparam ss_4__I_0_319_i9_2_lut_rep_438_3_lut_4_lut.init = 16'hfdff;
    LUT4 equal_114_i9_2_lut_rep_431_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21894), 
         .D(n22379), .Z(n21851)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(175[9:17])
    defparam equal_114_i9_2_lut_rep_431_3_lut_4_lut.init = 16'hfdff;
    LUT4 i13584_2_lut (.A(addOut[12]), .B(n22388), .Z(backOut1_28__N_1445[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13584_2_lut.init = 16'h2222;
    LUT4 i3426_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m2[18]), .Z(n5723)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3426_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3428_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m2[19]), .Z(n5725)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3428_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i29_4_lut (.A(backOut2_c[28]), .B(backOut3_c[28]), .C(n21851), 
         .D(n9), .Z(n558[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i29_4_lut.init = 16'h0aca;
    LUT4 mux_198_i4_3_lut_4_lut_3_lut (.A(n1145[15]), .B(n30_adj_1851), 
         .C(n2153[3]), .Z(n1258[3])) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(326[7:42])
    defparam mux_198_i4_3_lut_4_lut_3_lut.init = 16'ha2a2;
    CCU2D add_179_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[13]), .B1(n19130), .C1(n19131), .D1(Out0[28]), .COUT(n18682), 
          .S1(n1145[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(314[17:21])
    defparam add_179_1.INIT0 = 16'hF000;
    defparam add_179_1.INIT1 = 16'h56aa;
    defparam add_179_1.INJECT1_0 = "NO";
    defparam add_179_1.INJECT1_1 = "NO";
    CCU2D add_1180_23 (.A0(n5178), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18681), 
          .S0(n2245[21]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_23.INIT0 = 16'hf555;
    defparam add_1180_23.INIT1 = 16'h0000;
    defparam add_1180_23.INJECT1_0 = "NO";
    defparam add_1180_23.INJECT1_1 = "NO";
    CCU2D add_16131_21 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18878), .S1(n42));
    defparam add_16131_21.INIT0 = 16'h5555;
    defparam add_16131_21.INIT1 = 16'h0000;
    defparam add_16131_21.INJECT1_0 = "NO";
    defparam add_16131_21.INJECT1_1 = "NO";
    CCU2D add_16131_19 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18877), .COUT(n18878));
    defparam add_16131_19.INIT0 = 16'hf555;
    defparam add_16131_19.INIT1 = 16'hf555;
    defparam add_16131_19.INJECT1_0 = "NO";
    defparam add_16131_19.INJECT1_1 = "NO";
    LUT4 i3432_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m2[20]), .Z(n5729)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3432_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i21_4_lut (.A(backOut2_c[20]), .B(backOut3_c[20]), .C(n21851), 
         .D(n9), .Z(n558[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i21_4_lut.init = 16'h0aca;
    CCU2D add_1180_21 (.A0(n5176), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5178), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18680), 
          .COUT(n18681), .S0(n2245[19]), .S1(n2245[20]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_21.INIT0 = 16'hf555;
    defparam add_1180_21.INIT1 = 16'hf555;
    defparam add_1180_21.INJECT1_0 = "NO";
    defparam add_1180_21.INJECT1_1 = "NO";
    LUT4 i13583_2_lut (.A(addOut[11]), .B(n22388), .Z(backOut1_28__N_1445[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13583_2_lut.init = 16'h2222;
    CCU2D add_16131_17 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18876), .COUT(n18877));
    defparam add_16131_17.INIT0 = 16'hf555;
    defparam add_16131_17.INIT1 = 16'hf555;
    defparam add_16131_17.INJECT1_0 = "NO";
    defparam add_16131_17.INJECT1_1 = "NO";
    LUT4 i13582_2_lut (.A(addOut[10]), .B(n22388), .Z(backOut1_28__N_1445[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13582_2_lut.init = 16'h2222;
    CCU2D add_1180_19 (.A0(n5172), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5174), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18679), 
          .COUT(n18680), .S0(n2245[17]), .S1(n2245[18]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_19.INIT0 = 16'hf555;
    defparam add_1180_19.INIT1 = 16'hf555;
    defparam add_1180_19.INJECT1_0 = "NO";
    defparam add_1180_19.INJECT1_1 = "NO";
    LUT4 i13593_2_lut (.A(addOut[9]), .B(n22388), .Z(backOut2_28__N_1474[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13593_2_lut.init = 16'h2222;
    CCU2D add_16131_15 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18875), .COUT(n18876));
    defparam add_16131_15.INIT0 = 16'hf555;
    defparam add_16131_15.INIT1 = 16'hf555;
    defparam add_16131_15.INJECT1_0 = "NO";
    defparam add_16131_15.INJECT1_1 = "NO";
    LUT4 i2960_3_lut_4_lut (.A(n21824), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m2[0]), .Z(n5254)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i2960_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i12_4_lut (.A(backOut2_c[11]), .B(backOut3_c[11]), .C(n21851), 
         .D(n9), .Z(n558[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i12_4_lut.init = 16'h0aca;
    LUT4 i13592_2_lut (.A(addOut[8]), .B(n22388), .Z(backOut2_28__N_1474[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13592_2_lut.init = 16'h2222;
    LUT4 i13611_2_lut (.A(addOut[7]), .B(n22388), .Z(Out0_28__N_853[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13611_2_lut.init = 16'h2222;
    LUT4 mux_198_i6_3_lut_4_lut_3_lut (.A(n1145[15]), .B(n30_adj_1851), 
         .C(n2153[5]), .Z(n1258[5])) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(326[7:42])
    defparam mux_198_i6_3_lut_4_lut_3_lut.init = 16'ha2a2;
    LUT4 mux_135_i22_4_lut (.A(backOut2_c[21]), .B(backOut3_c[21]), .C(n21851), 
         .D(n9), .Z(n558[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i22_4_lut.init = 16'h0aca;
    LUT4 mux_198_i8_3_lut_4_lut_3_lut (.A(n1145[15]), .B(n30_adj_1851), 
         .C(n2153[7]), .Z(n1258[7])) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(326[7:42])
    defparam mux_198_i8_3_lut_4_lut_3_lut.init = 16'ha2a2;
    CCU2D add_16131_13 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18874), .COUT(n18875));
    defparam add_16131_13.INIT0 = 16'hf555;
    defparam add_16131_13.INIT1 = 16'hf555;
    defparam add_16131_13.INJECT1_0 = "NO";
    defparam add_16131_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_106 (.A(ss[1]), .B(n20184), .C(n22388), .D(n20055), 
         .Z(clk_N_683_enable_324)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_106.init = 16'hc4c0;
    LUT4 mux_135_i13_4_lut (.A(backOut2_c[12]), .B(backOut3_c[12]), .C(n21851), 
         .D(n9), .Z(n558[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i13_4_lut.init = 16'h0aca;
    CCU2D add_16122_21 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18991), .S1(n49));
    defparam add_16122_21.INIT0 = 16'h5555;
    defparam add_16122_21.INIT1 = 16'h0000;
    defparam add_16122_21.INJECT1_0 = "NO";
    defparam add_16122_21.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_107 (.A(ss[1]), .B(n20184), .C(n22388), .D(n20055), 
         .Z(clk_N_683_enable_352)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_107.init = 16'hc8c0;
    CCU2D add_16122_19 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18990), .COUT(n18991));
    defparam add_16122_19.INIT0 = 16'hf555;
    defparam add_16122_19.INIT1 = 16'hf555;
    defparam add_16122_19.INJECT1_0 = "NO";
    defparam add_16122_19.INJECT1_1 = "NO";
    LUT4 mux_135_i14_4_lut (.A(backOut2_c[13]), .B(backOut3_c[13]), .C(n21851), 
         .D(n9), .Z(n558[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i14_4_lut.init = 16'h0aca;
    LUT4 mux_135_i23_4_lut (.A(backOut2_c[22]), .B(backOut3_c[22]), .C(n21851), 
         .D(n9), .Z(n558[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i23_4_lut.init = 16'h0aca;
    LUT4 i13581_2_lut (.A(addOut[6]), .B(n22388), .Z(backOut1_28__N_1445[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13581_2_lut.init = 16'h2222;
    LUT4 mux_135_i24_4_lut (.A(backOut2_c[23]), .B(backOut3_c[23]), .C(n21851), 
         .D(n9), .Z(n558[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i24_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_108 (.A(n21886), .B(n20184), .C(n22388), .D(n21924), 
         .Z(clk_N_683_enable_72)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_108.init = 16'hc4c0;
    CCU2D add_1180_17 (.A0(n5168), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5170), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18678), 
          .COUT(n18679), .S0(n2245[15]), .S1(n2245[16]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_17.INIT0 = 16'hf555;
    defparam add_1180_17.INIT1 = 16'hf555;
    defparam add_1180_17.INJECT1_0 = "NO";
    defparam add_1180_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_109 (.A(n22388), .B(addOut[5]), .Z(backOut2_28__N_1474[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_adj_109.init = 16'h4444;
    CCU2D add_16122_17 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18989), .COUT(n18990));
    defparam add_16122_17.INIT0 = 16'hf555;
    defparam add_16122_17.INIT1 = 16'hf555;
    defparam add_16122_17.INJECT1_0 = "NO";
    defparam add_16122_17.INJECT1_1 = "NO";
    CCU2D add_16122_15 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18988), .COUT(n18989));
    defparam add_16122_15.INIT0 = 16'hf555;
    defparam add_16122_15.INIT1 = 16'hf555;
    defparam add_16122_15.INJECT1_0 = "NO";
    defparam add_16122_15.INJECT1_1 = "NO";
    LUT4 mux_135_i15_4_lut (.A(backOut2_c[14]), .B(backOut3_c[14]), .C(n21851), 
         .D(n9), .Z(n558[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i15_4_lut.init = 16'h0aca;
    CCU2D add_16122_13 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18987), .COUT(n18988));
    defparam add_16122_13.INIT0 = 16'hf555;
    defparam add_16122_13.INIT1 = 16'hf555;
    defparam add_16122_13.INJECT1_0 = "NO";
    defparam add_16122_13.INJECT1_1 = "NO";
    CCU2D add_16122_11 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18986), .COUT(n18987));
    defparam add_16122_11.INIT0 = 16'hf555;
    defparam add_16122_11.INIT1 = 16'hf555;
    defparam add_16122_11.INJECT1_0 = "NO";
    defparam add_16122_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_110 (.A(n22388), .B(addOut[4]), .Z(backOut1_28__N_1445[4])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_adj_110.init = 16'h4444;
    CCU2D add_16122_9 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18985), .COUT(n18986));
    defparam add_16122_9.INIT0 = 16'hf555;
    defparam add_16122_9.INIT1 = 16'hf555;
    defparam add_16122_9.INJECT1_0 = "NO";
    defparam add_16122_9.INJECT1_1 = "NO";
    LUT4 mux_135_i16_4_lut (.A(backOut2_c[15]), .B(backOut3_c[15]), .C(n21851), 
         .D(n9), .Z(n558[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(184[17] 191[27])
    defparam mux_135_i16_4_lut.init = 16'h0aca;
    CCU2D add_16131_11 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18873), .COUT(n18874));
    defparam add_16131_11.INIT0 = 16'hf555;
    defparam add_16131_11.INIT1 = 16'hf555;
    defparam add_16131_11.INJECT1_0 = "NO";
    defparam add_16131_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_111 (.A(n22388), .B(addOut[3]), .Z(backOut2_28__N_1474[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_adj_111.init = 16'h4444;
    CCU2D add_16131_9 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18872), .COUT(n18873));
    defparam add_16131_9.INIT0 = 16'hf555;
    defparam add_16131_9.INIT1 = 16'hf555;
    defparam add_16131_9.INJECT1_0 = "NO";
    defparam add_16131_9.INJECT1_1 = "NO";
    CCU2D add_16122_7 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18984), .COUT(n18985));
    defparam add_16122_7.INIT0 = 16'hf555;
    defparam add_16122_7.INIT1 = 16'hf555;
    defparam add_16122_7.INJECT1_0 = "NO";
    defparam add_16122_7.INJECT1_1 = "NO";
    CCU2D add_1177_11 (.A0(n1208[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18780), 
          .S0(n2189[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(351[20:29])
    defparam add_1177_11.INIT0 = 16'hf555;
    defparam add_1177_11.INIT1 = 16'h0000;
    defparam add_1177_11.INJECT1_0 = "NO";
    defparam add_1177_11.INJECT1_1 = "NO";
    LUT4 mux_198_i7_3_lut_4_lut_3_lut (.A(n1145[15]), .B(n30_adj_1851), 
         .C(n2153[6]), .Z(n1258[6])) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(326[7:42])
    defparam mux_198_i7_3_lut_4_lut_3_lut.init = 16'ha2a2;
    CCU2D add_16122_5 (.A0(speed_set_m3[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18983), .COUT(n18984));
    defparam add_16122_5.INIT0 = 16'hf555;
    defparam add_16122_5.INIT1 = 16'hf555;
    defparam add_16122_5.INJECT1_0 = "NO";
    defparam add_16122_5.INJECT1_1 = "NO";
    CCU2D add_16131_7 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18871), .COUT(n18872));
    defparam add_16131_7.INIT0 = 16'hf555;
    defparam add_16131_7.INIT1 = 16'hf555;
    defparam add_16131_7.INJECT1_0 = "NO";
    defparam add_16131_7.INJECT1_1 = "NO";
    CCU2D add_16122_3 (.A0(speed_set_m3[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18982), .COUT(n18983));
    defparam add_16122_3.INIT0 = 16'hf555;
    defparam add_16122_3.INIT1 = 16'hf555;
    defparam add_16122_3.INJECT1_0 = "NO";
    defparam add_16122_3.INJECT1_1 = "NO";
    CCU2D add_16122_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[0]), .B1(speed_set_m3[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18982));
    defparam add_16122_1.INIT0 = 16'hF000;
    defparam add_16122_1.INIT1 = 16'ha666;
    defparam add_16122_1.INJECT1_0 = "NO";
    defparam add_16122_1.INJECT1_1 = "NO";
    CCU2D add_16123_21 (.A0(speed_set_m1[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18981), .S1(n35));
    defparam add_16123_21.INIT0 = 16'h5555;
    defparam add_16123_21.INIT1 = 16'h0000;
    defparam add_16123_21.INJECT1_0 = "NO";
    defparam add_16123_21.INJECT1_1 = "NO";
    CCU2D add_16123_19 (.A0(speed_set_m1[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18980), .COUT(n18981));
    defparam add_16123_19.INIT0 = 16'hf555;
    defparam add_16123_19.INIT1 = 16'hf555;
    defparam add_16123_19.INJECT1_0 = "NO";
    defparam add_16123_19.INJECT1_1 = "NO";
    CCU2D add_1180_15 (.A0(n5164), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5166), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18677), 
          .COUT(n18678), .S0(n2245[13]), .S1(n2245[14]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_15.INIT0 = 16'hf555;
    defparam add_1180_15.INIT1 = 16'hf555;
    defparam add_1180_15.INJECT1_0 = "NO";
    defparam add_1180_15.INJECT1_1 = "NO";
    CCU2D add_16123_17 (.A0(speed_set_m1[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18979), .COUT(n18980));
    defparam add_16123_17.INIT0 = 16'hf555;
    defparam add_16123_17.INIT1 = 16'hf555;
    defparam add_16123_17.INJECT1_0 = "NO";
    defparam add_16123_17.INJECT1_1 = "NO";
    CCU2D add_1177_9 (.A0(n1208[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18779), 
          .COUT(n18780), .S0(n2189[7]), .S1(n2189[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(351[20:29])
    defparam add_1177_9.INIT0 = 16'hf555;
    defparam add_1177_9.INIT1 = 16'hf555;
    defparam add_1177_9.INJECT1_0 = "NO";
    defparam add_1177_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_112 (.A(n22388), .B(addOut[2]), .Z(backOut3_28__N_1503[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_adj_112.init = 16'h4444;
    LUT4 i1_2_lut_adj_113 (.A(n22388), .B(addOut[1]), .Z(backOut2_28__N_1474[1])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_adj_113.init = 16'h4444;
    PFUMX mux_1194_i21 (.BLUT(n5130), .ALUT(n5088), .C0(n2437), .Z(n5178));
    CCU2D add_16123_15 (.A0(speed_set_m1[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18978), .COUT(n18979));
    defparam add_16123_15.INIT0 = 16'hf555;
    defparam add_16123_15.INIT1 = 16'hf555;
    defparam add_16123_15.INJECT1_0 = "NO";
    defparam add_16123_15.INJECT1_1 = "NO";
    CCU2D add_16123_13 (.A0(speed_set_m1[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18977), .COUT(n18978));
    defparam add_16123_13.INIT0 = 16'hf555;
    defparam add_16123_13.INIT1 = 16'hf555;
    defparam add_16123_13.INJECT1_0 = "NO";
    defparam add_16123_13.INJECT1_1 = "NO";
    CCU2D add_16123_11 (.A0(speed_set_m1[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18976), .COUT(n18977));
    defparam add_16123_11.INIT0 = 16'hf555;
    defparam add_16123_11.INIT1 = 16'hf555;
    defparam add_16123_11.INJECT1_0 = "NO";
    defparam add_16123_11.INJECT1_1 = "NO";
    PFUMX mux_1194_i20 (.BLUT(n5128), .ALUT(n5086), .C0(n2437), .Z(n5176));
    PFUMX mux_1194_i19 (.BLUT(n5126), .ALUT(n5084), .C0(n2437), .Z(n5174));
    PFUMX mux_1194_i18 (.BLUT(n5124), .ALUT(n5082), .C0(n2437), .Z(n5172));
    PFUMX mux_1194_i17 (.BLUT(n5122), .ALUT(n5080), .C0(n2437), .Z(n5170));
    PFUMX mux_1194_i16 (.BLUT(n5120), .ALUT(n5078), .C0(n2437), .Z(n5168));
    PFUMX mux_1194_i15 (.BLUT(n5118), .ALUT(n5076), .C0(n2437), .Z(n5166));
    PFUMX mux_1194_i14 (.BLUT(n5116), .ALUT(n5074), .C0(n2437), .Z(n5164));
    CCU2D add_16131_5 (.A0(speed_set_m2[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18870), .COUT(n18871));
    defparam add_16131_5.INIT0 = 16'hf555;
    defparam add_16131_5.INIT1 = 16'hf555;
    defparam add_16131_5.INJECT1_0 = "NO";
    defparam add_16131_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_114 (.A(n22388), .B(addOut[0]), .Z(backOut3_28__N_1503[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_adj_114.init = 16'h4444;
    PFUMX mux_1194_i13 (.BLUT(n5114), .ALUT(n5072), .C0(n2437), .Z(n5162));
    PFUMX mux_1194_i12 (.BLUT(n5112), .ALUT(n5070), .C0(n2437), .Z(n5160));
    LUT4 i10664_3_lut_4_lut (.A(n1145[15]), .B(n30_adj_1851), .C(n19129), 
         .D(clk_N_683_enable_392), .Z(n13080)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(326[7:42])
    defparam i10664_3_lut_4_lut.init = 16'hf700;
    CCU2D add_16123_9 (.A0(speed_set_m1[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18975), .COUT(n18976));
    defparam add_16123_9.INIT0 = 16'hf555;
    defparam add_16123_9.INIT1 = 16'hf555;
    defparam add_16123_9.INJECT1_0 = "NO";
    defparam add_16123_9.INJECT1_1 = "NO";
    PFUMX mux_1194_i11 (.BLUT(n5110), .ALUT(n5068), .C0(n2437), .Z(n5158));
    PFUMX mux_1194_i10 (.BLUT(n5108), .ALUT(n5066), .C0(n2437), .Z(n5156));
    CCU2D add_16123_7 (.A0(speed_set_m1[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18974), .COUT(n18975));
    defparam add_16123_7.INIT0 = 16'hf555;
    defparam add_16123_7.INIT1 = 16'hf555;
    defparam add_16123_7.INJECT1_0 = "NO";
    defparam add_16123_7.INJECT1_1 = "NO";
    CCU2D add_16131_3 (.A0(speed_set_m2[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18869), .COUT(n18870));
    defparam add_16131_3.INIT0 = 16'hf555;
    defparam add_16131_3.INIT1 = 16'hf555;
    defparam add_16131_3.INJECT1_0 = "NO";
    defparam add_16131_3.INJECT1_1 = "NO";
    CCU2D add_16123_5 (.A0(speed_set_m1[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18973), .COUT(n18974));
    defparam add_16123_5.INIT0 = 16'hf555;
    defparam add_16123_5.INIT1 = 16'hf555;
    defparam add_16123_5.INJECT1_0 = "NO";
    defparam add_16123_5.INJECT1_1 = "NO";
    CCU2D add_16123_3 (.A0(speed_set_m1[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18972), .COUT(n18973));
    defparam add_16123_3.INIT0 = 16'hf555;
    defparam add_16123_3.INIT1 = 16'hf555;
    defparam add_16123_3.INJECT1_0 = "NO";
    defparam add_16123_3.INJECT1_1 = "NO";
    PFUMX mux_1194_i9 (.BLUT(n5106), .ALUT(n5064), .C0(n2437), .Z(n5154));
    PFUMX mux_1194_i8 (.BLUT(n5104), .ALUT(n5062), .C0(n2437), .Z(n5152));
    PFUMX mux_1194_i7 (.BLUT(n5102), .ALUT(n5060), .C0(n2437), .Z(n5150));
    PFUMX mux_1194_i6 (.BLUT(n5100), .ALUT(n5058), .C0(n2437), .Z(n5148));
    PFUMX mux_1194_i5 (.BLUT(n5098), .ALUT(n5056), .C0(n2437), .Z(n5146));
    PFUMX mux_1194_i4 (.BLUT(n5096), .ALUT(n5054), .C0(n2437), .Z(n5144));
    PFUMX mux_1194_i3 (.BLUT(n5094), .ALUT(n5052), .C0(n2437), .Z(n5142));
    PFUMX mux_1194_i2 (.BLUT(n5092), .ALUT(n5050), .C0(n2437), .Z(n5140));
    PFUMX mux_1194_i1 (.BLUT(n5048), .ALUT(n5046), .C0(n2437), .Z(n5138));
    PFUMX i3393 (.BLUT(n2485[1]), .ALUT(n5689), .C0(n21815), .Z(n5690));
    PFUMX i3395 (.BLUT(n2485[2]), .ALUT(n5691), .C0(n21815), .Z(n5692));
    LUT4 i3434_2_lut_rep_470 (.A(n22388), .B(n22383), .Z(clk_N_683_enable_392)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i3434_2_lut_rep_470.init = 16'h8888;
    CCU2D add_16123_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[0]), .B1(speed_set_m1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18972));
    defparam add_16123_1.INIT0 = 16'hF000;
    defparam add_16123_1.INIT1 = 16'ha666;
    defparam add_16123_1.INJECT1_0 = "NO";
    defparam add_16123_1.INJECT1_1 = "NO";
    CCU2D add_16131_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[0]), .B1(speed_set_m2[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18869));
    defparam add_16131_1.INIT0 = 16'hF000;
    defparam add_16131_1.INIT1 = 16'ha666;
    defparam add_16131_1.INJECT1_0 = "NO";
    defparam add_16131_1.INJECT1_1 = "NO";
    LUT4 i10807_2_lut_3_lut_4_lut (.A(n22388), .B(n22383), .C(n21922), 
         .D(n21923), .Z(n13082)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i10807_2_lut_3_lut_4_lut.init = 16'h8880;
    PFUMX i3397 (.BLUT(n2485[3]), .ALUT(n5693), .C0(n21815), .Z(n5694));
    PFUMX i3399 (.BLUT(n2485[4]), .ALUT(n5695), .C0(n21815), .Z(n5696));
    PFUMX i3401 (.BLUT(n2485[5]), .ALUT(n5697), .C0(n21815), .Z(n5698));
    PFUMX i3403 (.BLUT(n2485[6]), .ALUT(n5699), .C0(n21815), .Z(n5700));
    CCU2D add_16121_21 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18868), .S1(n56));
    defparam add_16121_21.INIT0 = 16'h5555;
    defparam add_16121_21.INIT1 = 16'h0000;
    defparam add_16121_21.INJECT1_0 = "NO";
    defparam add_16121_21.INJECT1_1 = "NO";
    PFUMX i3405 (.BLUT(n2485[7]), .ALUT(n5701), .C0(n21815), .Z(n5702));
    PFUMX i3407 (.BLUT(n2485[8]), .ALUT(n5703), .C0(n21815), .Z(n5704));
    PFUMX i3409 (.BLUT(n2485[9]), .ALUT(n5705), .C0(n21815), .Z(n5706));
    PFUMX i3411 (.BLUT(n2485[10]), .ALUT(n5707), .C0(n21815), .Z(n5708));
    CCU2D add_16121_19 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18867), .COUT(n18868));
    defparam add_16121_19.INIT0 = 16'hf555;
    defparam add_16121_19.INIT1 = 16'hf555;
    defparam add_16121_19.INJECT1_0 = "NO";
    defparam add_16121_19.INJECT1_1 = "NO";
    LUT4 i13274_2_lut_rep_472 (.A(ss[0]), .B(ss[1]), .Z(n21892)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i13274_2_lut_rep_472.init = 16'h8888;
    PFUMX i3413 (.BLUT(n2485[11]), .ALUT(n5709), .C0(n21815), .Z(n5710));
    CCU2D add_16121_17 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18866), .COUT(n18867));
    defparam add_16121_17.INIT0 = 16'hf555;
    defparam add_16121_17.INIT1 = 16'hf555;
    defparam add_16121_17.INJECT1_0 = "NO";
    defparam add_16121_17.INJECT1_1 = "NO";
    PFUMX i3415 (.BLUT(n2485[12]), .ALUT(n5711), .C0(n21815), .Z(n5712));
    PFUMX i3417 (.BLUT(n2485[13]), .ALUT(n5713), .C0(n21815), .Z(n5714));
    PFUMX i3419 (.BLUT(n2485[14]), .ALUT(n5715), .C0(n21815), .Z(n5716));
    PFUMX i3421 (.BLUT(n2485[15]), .ALUT(n5717), .C0(n21815), .Z(n5718));
    CCU2D add_16121_15 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18865), .COUT(n18866));
    defparam add_16121_15.INIT0 = 16'hf555;
    defparam add_16121_15.INIT1 = 16'hf555;
    defparam add_16121_15.INJECT1_0 = "NO";
    defparam add_16121_15.INJECT1_1 = "NO";
    PFUMX i3423 (.BLUT(n2485[16]), .ALUT(n5719), .C0(n21815), .Z(n5720));
    PFUMX i3425 (.BLUT(n2485[17]), .ALUT(n5721), .C0(n21815), .Z(n5722));
    PFUMX i3427 (.BLUT(n2485[18]), .ALUT(n5723), .C0(n21815), .Z(n5724));
    CCU2D add_16121_13 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18864), .COUT(n18865));
    defparam add_16121_13.INIT0 = 16'hf555;
    defparam add_16121_13.INIT1 = 16'hf555;
    defparam add_16121_13.INJECT1_0 = "NO";
    defparam add_16121_13.INJECT1_1 = "NO";
    CCU2D add_16121_11 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18863), .COUT(n18864));
    defparam add_16121_11.INIT0 = 16'hf555;
    defparam add_16121_11.INIT1 = 16'hf555;
    defparam add_16121_11.INJECT1_0 = "NO";
    defparam add_16121_11.INJECT1_1 = "NO";
    PFUMX i3429 (.BLUT(n2485[19]), .ALUT(n5725), .C0(n21815), .Z(n5726));
    PFUMX i3433 (.BLUT(n2485[20]), .ALUT(n5729), .C0(n21815), .Z(n5730));
    LUT4 i1_2_lut_rep_430_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21893), 
         .D(n22379), .Z(n21850)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_430_3_lut_4_lut.init = 16'hfff7;
    PFUMX i2961 (.BLUT(n2485[0]), .ALUT(n5254), .C0(n21815), .Z(n5255));
    CCU2D add_16121_9 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18862), .COUT(n18863));
    defparam add_16121_9.INIT0 = 16'hf555;
    defparam add_16121_9.INIT1 = 16'hf555;
    defparam add_16121_9.INJECT1_0 = "NO";
    defparam add_16121_9.INJECT1_1 = "NO";
    CCU2D add_16121_7 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18861), .COUT(n18862));
    defparam add_16121_7.INIT0 = 16'hf555;
    defparam add_16121_7.INIT1 = 16'hf555;
    defparam add_16121_7.INJECT1_0 = "NO";
    defparam add_16121_7.INJECT1_1 = "NO";
    LUT4 equal_110_i9_2_lut_rep_428_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21894), 
         .D(ss[2]), .Z(n21848)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam equal_110_i9_2_lut_rep_428_3_lut_4_lut.init = 16'hfff7;
    L6MUX21 addIn2_28__I_29_i29 (.D0(n618[28]), .D1(addIn2_28__N_1337[28]), 
            .SD(n20537), .Z(addIn2_28__N_1207[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i28 (.D0(n618[27]), .D1(addIn2_28__N_1337[27]), 
            .SD(n20537), .Z(addIn2_28__N_1207[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i27 (.D0(n618[26]), .D1(addIn2_28__N_1337[26]), 
            .SD(n20537), .Z(addIn2_28__N_1207[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i26 (.D0(n618[25]), .D1(addIn2_28__N_1337[25]), 
            .SD(n20537), .Z(addIn2_28__N_1207[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i25 (.D0(n618[24]), .D1(addIn2_28__N_1337[24]), 
            .SD(n20537), .Z(addIn2_28__N_1207[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i24 (.D0(n618[23]), .D1(addIn2_28__N_1337[23]), 
            .SD(n20537), .Z(addIn2_28__N_1207[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i23 (.D0(n618[22]), .D1(addIn2_28__N_1337[22]), 
            .SD(n20537), .Z(addIn2_28__N_1207[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 ss_4__I_0_321_i9_2_lut_rep_442_3_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21893), .D(ss[2]), .Z(n21862)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam ss_4__I_0_321_i9_2_lut_rep_442_3_lut_4_lut.init = 16'hf7ff;
    L6MUX21 addIn2_28__I_29_i22 (.D0(n618[21]), .D1(addIn2_28__N_1337[21]), 
            .SD(n20537), .Z(addIn2_28__N_1207[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i21 (.D0(n618[20]), .D1(addIn2_28__N_1337[20]), 
            .SD(n20537), .Z(addIn2_28__N_1207[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i20 (.D0(n618[19]), .D1(addIn2_28__N_1337[19]), 
            .SD(n20537), .Z(addIn2_28__N_1207[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_16121_5 (.A0(speed_set_m4[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18860), .COUT(n18861));
    defparam add_16121_5.INIT0 = 16'hf555;
    defparam add_16121_5.INIT1 = 16'hf555;
    defparam add_16121_5.INJECT1_0 = "NO";
    defparam add_16121_5.INJECT1_1 = "NO";
    CCU2D add_16121_3 (.A0(speed_set_m4[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18859), .COUT(n18860));
    defparam add_16121_3.INIT0 = 16'hf555;
    defparam add_16121_3.INIT1 = 16'hf555;
    defparam add_16121_3.INJECT1_0 = "NO";
    defparam add_16121_3.INJECT1_1 = "NO";
    L6MUX21 addIn2_28__I_29_i19 (.D0(n618[18]), .D1(addIn2_28__N_1337[18]), 
            .SD(n20537), .Z(addIn2_28__N_1207[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i7790_2_lut_3_lut (.A(ss[0]), .B(ss[1]), .C(ss[2]), .Z(n14_c)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i7790_2_lut_3_lut.init = 16'h7878;
    L6MUX21 addIn2_28__I_29_i18 (.D0(n618[17]), .D1(addIn2_28__N_1337[17]), 
            .SD(n20537), .Z(addIn2_28__N_1207[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i9 (.D0(n618[8]), .D1(addIn2_28__N_1337[8]), 
            .SD(n20537), .Z(addIn2_28__N_1207[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i7_4_lut_adj_115 (.A(Out1[3]), .B(n14_adj_1858), .C(n10_adj_1859), 
         .D(Out1[4]), .Z(n19086)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam i7_4_lut_adj_115.init = 16'hfffe;
    L6MUX21 addIn2_28__I_29_i7 (.D0(n618[6]), .D1(addIn2_28__N_1337[6]), 
            .SD(n20537), .Z(addIn2_28__N_1207[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_198_i10_3_lut_4_lut_3_lut (.A(n1145[15]), .B(n30_adj_1851), 
         .C(n2153[9]), .Z(n1258[9])) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(326[7:42])
    defparam mux_198_i10_3_lut_4_lut_3_lut.init = 16'ha2a2;
    L6MUX21 addIn2_28__I_29_i8 (.D0(n618[7]), .D1(addIn2_28__N_1337[7]), 
            .SD(n20537), .Z(addIn2_28__N_1207[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i10 (.D0(n618[9]), .D1(addIn2_28__N_1337[9]), 
            .SD(n20537), .Z(addIn2_28__N_1207[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i11 (.D0(n618[10]), .D1(addIn2_28__N_1337[10]), 
            .SD(n20537), .Z(addIn2_28__N_1207[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i12 (.D0(n618[11]), .D1(addIn2_28__N_1337[11]), 
            .SD(n20537), .Z(addIn2_28__N_1207[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i13 (.D0(n618[12]), .D1(addIn2_28__N_1337[12]), 
            .SD(n20537), .Z(addIn2_28__N_1207[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i14 (.D0(n618[13]), .D1(addIn2_28__N_1337[13]), 
            .SD(n20537), .Z(addIn2_28__N_1207[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i6_4_lut_adj_116 (.A(Out1[11]), .B(Out1[7]), .C(Out1[2]), .D(Out1[10]), 
         .Z(n14_adj_1858)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam i6_4_lut_adj_116.init = 16'hfffe;
    L6MUX21 addIn2_28__I_29_i15 (.D0(n618[14]), .D1(addIn2_28__N_1337[14]), 
            .SD(n20537), .Z(addIn2_28__N_1207[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i16 (.D0(n618[15]), .D1(addIn2_28__N_1337[15]), 
            .SD(n20537), .Z(addIn2_28__N_1207[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    L6MUX21 addIn2_28__I_29_i17 (.D0(n618[16]), .D1(addIn2_28__N_1337[16]), 
            .SD(n20537), .Z(addIn2_28__N_1207[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_1802_i4 (.BLUT(n3691[3]), .ALUT(subIn2_24__N_1114[3]), .C0(n20582), 
          .Z(subIn2[3]));
    LUT4 i2_2_lut_adj_117 (.A(Out1[9]), .B(Out1[1]), .Z(n10_adj_1859)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam i2_2_lut_adj_117.init = 16'heeee;
    CCU2D add_16121_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[0]), .B1(speed_set_m4[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18859));
    defparam add_16121_1.INIT0 = 16'hF000;
    defparam add_16121_1.INIT1 = 16'ha666;
    defparam add_16121_1.INJECT1_0 = "NO";
    defparam add_16121_1.INJECT1_1 = "NO";
    PFUMX mux_1802_i8 (.BLUT(n3691[7]), .ALUT(subIn2_24__N_1114[7]), .C0(n20582), 
          .Z(subIn2[7]));
    PFUMX mux_1802_i9 (.BLUT(n3691[8]), .ALUT(subIn2_24__N_1114[8]), .C0(n20582), 
          .Z(subIn2[8]));
    CCU2D sub_17_rep_3_add_2_23 (.A0(n21816), .B0(n16318), .C0(n57), .D0(n5730), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18858), 
          .S0(n4208));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_23.INIT0 = 16'h04ff;
    defparam sub_17_rep_3_add_2_23.INIT1 = 16'h0000;
    defparam sub_17_rep_3_add_2_23.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_23.INJECT1_1 = "NO";
    PFUMX mux_1802_i10 (.BLUT(n3691[9]), .ALUT(subIn2_24__N_1114[9]), .C0(n20582), 
          .Z(subIn2[9]));
    LUT4 i13201_2_lut_rep_473 (.A(n22388), .B(ss[3]), .Z(n21893)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13201_2_lut_rep_473.init = 16'heeee;
    LUT4 i4_4_lut_adj_118 (.A(Out1[5]), .B(Out1[6]), .C(Out1[0]), .D(n6_adj_1860), 
         .Z(n19087)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam i4_4_lut_adj_118.init = 16'hfffe;
    LUT4 ss_4__I_0_314_i6_2_lut (.A(ss[0]), .B(ss[1]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(165[9:16])
    defparam ss_4__I_0_314_i6_2_lut.init = 16'heeee;
    PFUMX mux_1802_i13 (.BLUT(n3691[12]), .ALUT(subIn2_24__N_1114[12]), 
          .C0(n20582), .Z(subIn2[12]));
    LUT4 i1_2_lut_adj_119 (.A(Out1[8]), .B(Out1[12]), .Z(n6_adj_1860)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam i1_2_lut_adj_119.init = 16'heeee;
    LUT4 i1_2_lut_rep_447_3_lut (.A(n22388), .B(ss[3]), .C(n22379), .Z(n21867)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_447_3_lut.init = 16'hfefe;
    CCU2D sub_17_rep_3_add_2_21 (.A0(n7), .B0(n16318), .C0(n16214), .D0(n5726), 
          .A1(n21816), .B1(n16318), .C1(n57), .D1(n5730), .CIN(n18857), 
          .COUT(n18858), .S0(n4210), .S1(n4209));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_21.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_21.INIT1 = 16'h04ff;
    defparam sub_17_rep_3_add_2_21.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_21.INJECT1_1 = "NO";
    CCU2D add_1177_7 (.A0(n1208[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18778), 
          .COUT(n18779), .S0(n2189[5]), .S1(n2189[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(351[20:29])
    defparam add_1177_7.INIT0 = 16'hf555;
    defparam add_1177_7.INIT1 = 16'hf555;
    defparam add_1177_7.INJECT1_0 = "NO";
    defparam add_1177_7.INJECT1_1 = "NO";
    CCU2D add_1177_5 (.A0(n1208[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18777), 
          .COUT(n18778), .S0(n2189[3]), .S1(n2189[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(351[20:29])
    defparam add_1177_5.INIT0 = 16'hf555;
    defparam add_1177_5.INIT1 = 16'hf555;
    defparam add_1177_5.INJECT1_0 = "NO";
    defparam add_1177_5.INJECT1_1 = "NO";
    CCU2D sub_17_rep_3_add_2_19 (.A0(subIn2[17]), .B0(n16318), .C0(n16214), 
          .D0(n5722), .A1(subIn2[18]), .B1(n16318), .C1(n16214), .D1(n5724), 
          .CIN(n18856), .COUT(n18857), .S0(n4212), .S1(n4211));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_19.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_19.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_19.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_17_rep_3_add_2_17 (.A0(subIn2[15]), .B0(n16318), .C0(n16214), 
          .D0(n5718), .A1(subIn2[16]), .B1(n16318), .C1(n16214), .D1(n5720), 
          .CIN(n18855), .COUT(n18856), .S0(n4214), .S1(n4213));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_17.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_17.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_17.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_449_3_lut (.A(n22388), .B(ss[3]), .C(n22379), .Z(n21869)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_449_3_lut.init = 16'hefef;
    PFUMX mux_1802_i2 (.BLUT(subIn2_24__N_1301[1]), .ALUT(subIn2_24__N_1114[1]), 
          .C0(n20586), .Z(subIn2[1]));
    CCU2D sub_17_rep_3_add_2_15 (.A0(subIn2[13]), .B0(n16318), .C0(n16214), 
          .D0(n5714), .A1(subIn2[14]), .B1(n16318), .C1(n16214), .D1(n5716), 
          .CIN(n18854), .COUT(n18855), .S0(n4216), .S1(n4215));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_15.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_15.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_15.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_15.INJECT1_1 = "NO";
    PFUMX mux_1802_i3 (.BLUT(subIn2_24__N_1301[2]), .ALUT(subIn2_24__N_1114[2]), 
          .C0(n20586), .Z(subIn2[2]));
    PFUMX mux_1802_i5 (.BLUT(subIn2_24__N_1301[4]), .ALUT(subIn2_24__N_1114[4]), 
          .C0(n20586), .Z(subIn2[4]));
    CCU2D sub_17_rep_3_add_2_13 (.A0(subIn2[11]), .B0(n16318), .C0(n16214), 
          .D0(n5710), .A1(subIn2[12]), .B1(n16318), .C1(n16214), .D1(n5712), 
          .CIN(n18853), .COUT(n18854), .S0(n4218), .S1(n4217));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_13.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_13.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_13.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_17_rep_3_add_2_11 (.A0(subIn2[9]), .B0(n16318), .C0(n16214), 
          .D0(n5706), .A1(subIn2[10]), .B1(n16318), .C1(n16214), .D1(n5708), 
          .CIN(n18852), .COUT(n18853), .S0(n4220), .S1(n4219));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_11.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_11.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_11.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_437_3_lut_4_lut (.A(n22388), .B(ss[3]), .C(n22379), 
         .D(n22375), .Z(n21857)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_437_3_lut_4_lut.init = 16'h1000;
    PFUMX mux_1802_i6 (.BLUT(subIn2_24__N_1301[5]), .ALUT(subIn2_24__N_1114[5]), 
          .C0(n20586), .Z(subIn2[5]));
    LUT4 mux_198_i9_3_lut_4_lut_3_lut (.A(n1145[15]), .B(n30_adj_1851), 
         .C(n2153[8]), .Z(n1258[8])) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(326[7:42])
    defparam mux_198_i9_3_lut_4_lut_3_lut.init = 16'ha2a2;
    PFUMX mux_1802_i7 (.BLUT(subIn2_24__N_1301[6]), .ALUT(subIn2_24__N_1114[6]), 
          .C0(n20586), .Z(subIn2[6]));
    LUT4 i1_2_lut_rep_474 (.A(n22388), .B(ss[3]), .Z(n21894)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(174[9:17])
    defparam i1_2_lut_rep_474.init = 16'hbbbb;
    CCU2D sub_17_rep_3_add_2_9 (.A0(subIn2[7]), .B0(n16318), .C0(n16214), 
          .D0(n5702), .A1(subIn2[8]), .B1(n16318), .C1(n16214), .D1(n5704), 
          .CIN(n18851), .COUT(n18852), .S0(n4222), .S1(n4221));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_9.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_9.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_9.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_448_3_lut (.A(n22388), .B(ss[3]), .C(n22379), .Z(n21868)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(174[9:17])
    defparam i1_2_lut_rep_448_3_lut.init = 16'hfbfb;
    CCU2D add_1177_3 (.A0(n1208[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18776), 
          .COUT(n18777), .S0(n2189[1]), .S1(n2189[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(351[20:29])
    defparam add_1177_3.INIT0 = 16'hf555;
    defparam add_1177_3.INIT1 = 16'hf555;
    defparam add_1177_3.INJECT1_0 = "NO";
    defparam add_1177_3.INJECT1_1 = "NO";
    PFUMX mux_1802_i11 (.BLUT(subIn2_24__N_1301[10]), .ALUT(subIn2_24__N_1114[10]), 
          .C0(n20586), .Z(subIn2[10]));
    CCU2D add_1177_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18776), 
          .S1(n2189[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(351[20:29])
    defparam add_1177_1.INIT0 = 16'hF000;
    defparam add_1177_1.INIT1 = 16'h0aaa;
    defparam add_1177_1.INJECT1_0 = "NO";
    defparam add_1177_1.INJECT1_1 = "NO";
    PFUMX mux_1802_i12 (.BLUT(subIn2_24__N_1301[11]), .ALUT(subIn2_24__N_1114[11]), 
          .C0(n20586), .Z(subIn2[11]));
    CCU2D sub_17_rep_3_add_2_7 (.A0(subIn2[5]), .B0(n16318), .C0(n16214), 
          .D0(n5698), .A1(subIn2[6]), .B1(n16318), .C1(n16214), .D1(n5700), 
          .CIN(n18850), .COUT(n18851), .S0(n4224), .S1(n4223));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_7.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_7.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_7.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_7.INJECT1_1 = "NO";
    PFUMX mux_1802_i14 (.BLUT(subIn2_24__N_1301[13]), .ALUT(subIn2_24__N_1114[13]), 
          .C0(n20586), .Z(subIn2[13]));
    CCU2D sub_17_rep_3_add_2_5 (.A0(subIn2[3]), .B0(n16318), .C0(n16214), 
          .D0(n5694), .A1(subIn2[4]), .B1(n16318), .C1(n16214), .D1(n5696), 
          .CIN(n18849), .COUT(n18850), .S0(n4226), .S1(n4225));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_5.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_5.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_5.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_5.INJECT1_1 = "NO";
    CCU2D add_1180_13 (.A0(n5160), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5162), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18676), 
          .COUT(n18677), .S0(n2245[11]), .S1(n2245[12]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_13.INIT0 = 16'hf555;
    defparam add_1180_13.INIT1 = 16'hf555;
    defparam add_1180_13.INJECT1_0 = "NO";
    defparam add_1180_13.INJECT1_1 = "NO";
    PFUMX mux_1802_i15 (.BLUT(subIn2_24__N_1301[14]), .ALUT(subIn2_24__N_1114[14]), 
          .C0(n20586), .Z(subIn2[14]));
    CCU2D sub_17_rep_3_add_2_3 (.A0(subIn2[1]), .B0(n16318), .C0(n16214), 
          .D0(n5690), .A1(subIn2[2]), .B1(n16318), .C1(n16214), .D1(n5692), 
          .CIN(n18848), .COUT(n18849), .S0(n4228), .S1(n4227));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_3.INIT0 = 16'ha655;
    defparam sub_17_rep_3_add_2_3.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_3.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_3.INJECT1_1 = "NO";
    LUT4 ss_4__I_0_317_i9_2_lut_rep_429_3_lut_4_lut (.A(n22388), .B(ss[3]), 
         .C(n21895), .D(n22379), .Z(n21849)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(174[9:17])
    defparam ss_4__I_0_317_i9_2_lut_rep_429_3_lut_4_lut.init = 16'hfffb;
    PFUMX mux_1802_i16 (.BLUT(subIn2_24__N_1301[15]), .ALUT(subIn2_24__N_1114[15]), 
          .C0(n20586), .Z(subIn2[15]));
    PFUMX mux_1802_i17 (.BLUT(subIn2_24__N_1301[16]), .ALUT(subIn2_24__N_1114[16]), 
          .C0(n20586), .Z(subIn2[16]));
    PFUMX mux_1802_i18 (.BLUT(subIn2_24__N_1301[17]), .ALUT(subIn2_24__N_1114[17]), 
          .C0(n20586), .Z(subIn2[17]));
    CCU2D sub_17_rep_3_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(subIn2[0]), .B1(n16318), .C1(n16214), .D1(n5255), 
          .COUT(n18848), .S1(n4229));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_3_add_2_1.INIT0 = 16'h0000;
    defparam sub_17_rep_3_add_2_1.INIT1 = 16'ha655;
    defparam sub_17_rep_3_add_2_1.INJECT1_0 = "NO";
    defparam sub_17_rep_3_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_463_3_lut (.A(n22388), .B(ss[3]), .C(ss[2]), .Z(n21883)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(174[9:17])
    defparam i1_2_lut_rep_463_3_lut.init = 16'hbfbf;
    CCU2D add_1176_11 (.A0(n1187[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18775), 
          .S0(n2177[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(343[20:29])
    defparam add_1176_11.INIT0 = 16'hf555;
    defparam add_1176_11.INIT1 = 16'h0000;
    defparam add_1176_11.INJECT1_0 = "NO";
    defparam add_1176_11.INJECT1_1 = "NO";
    CCU2D add_191_17 (.A0(Out3[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18713), 
          .S0(n1208[15]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_17.INIT0 = 16'h5aaa;
    defparam add_191_17.INIT1 = 16'h0000;
    defparam add_191_17.INJECT1_0 = "NO";
    defparam add_191_17.INJECT1_1 = "NO";
    LUT4 i10666_3_lut_4_lut (.A(n1166[15]), .B(n30_c), .C(n19129), .D(clk_N_683_enable_392), 
         .Z(n13089)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(334[7:42])
    defparam i10666_3_lut_4_lut.init = 16'hf700;
    CCU2D add_1176_9 (.A0(n1187[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18774), 
          .COUT(n18775), .S0(n2177[7]), .S1(n2177[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(343[20:29])
    defparam add_1176_9.INIT0 = 16'hf555;
    defparam add_1176_9.INIT1 = 16'hf555;
    defparam add_1176_9.INJECT1_0 = "NO";
    defparam add_1176_9.INJECT1_1 = "NO";
    LUT4 equal_133_i9_2_lut_3_lut_4_lut (.A(n22388), .B(ss[3]), .C(n21895), 
         .D(n22379), .Z(n9)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(174[9:17])
    defparam equal_133_i9_2_lut_3_lut_4_lut.init = 16'hfbff;
    CCU2D add_191_15 (.A0(Out3[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18712), 
          .COUT(n18713), .S0(n1208[13]), .S1(n1208[14]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_15.INIT0 = 16'h5aaa;
    defparam add_191_15.INIT1 = 16'h5aaa;
    defparam add_191_15.INJECT1_0 = "NO";
    defparam add_191_15.INJECT1_1 = "NO";
    CCU2D add_1180_11 (.A0(n5156), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5158), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18675), 
          .COUT(n18676), .S0(n2245[9]), .S1(n2245[10]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_11.INIT0 = 16'hf555;
    defparam add_1180_11.INIT1 = 16'hf555;
    defparam add_1180_11.INJECT1_0 = "NO";
    defparam add_1180_11.INJECT1_1 = "NO";
    LUT4 equal_133_i6_2_lut_rep_475 (.A(ss[0]), .B(ss[1]), .Z(n21895)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(192[19:27])
    defparam equal_133_i6_2_lut_rep_475.init = 16'hbbbb;
    LUT4 i13798_2_lut_rep_446_3_lut_2_lut (.A(ss[0]), .B(ss[1]), .Z(n21866)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(192[19:27])
    defparam i13798_2_lut_rep_446_3_lut_2_lut.init = 16'h9999;
    CCU2D add_1176_7 (.A0(n1187[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18773), 
          .COUT(n18774), .S0(n2177[5]), .S1(n2177[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(343[20:29])
    defparam add_1176_7.INIT0 = 16'hf555;
    defparam add_1176_7.INIT1 = 16'hf555;
    defparam add_1176_7.INJECT1_0 = "NO";
    defparam add_1176_7.INJECT1_1 = "NO";
    CCU2D add_191_13 (.A0(Out3[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18711), 
          .COUT(n18712), .S0(n1208[11]), .S1(n1208[12]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_13.INIT0 = 16'h5aaa;
    defparam add_191_13.INIT1 = 16'h5aaa;
    defparam add_191_13.INJECT1_0 = "NO";
    defparam add_191_13.INJECT1_1 = "NO";
    PFUMX mux_1802_i19 (.BLUT(subIn2_24__N_1301[18]), .ALUT(subIn2_24__N_1114[18]), 
          .C0(n20586), .Z(subIn2[18]));
    LUT4 mux_205_i7_3_lut_4_lut_3_lut (.A(n30_c), .B(n1166[15]), .C(n2165[6]), 
         .Z(n1302[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(334[25:42])
    defparam mux_205_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FD1S3IX ss_i2_rep_507 (.D(n14_c), .CK(clk_N_683), .CD(ss[4]), .Q(n22379));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam ss_i2_rep_507.GSR = "ENABLED";
    CCU2D add_1176_5 (.A0(n1187[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18772), 
          .COUT(n18773), .S0(n2177[3]), .S1(n2177[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(343[20:29])
    defparam add_1176_5.INIT0 = 16'hf555;
    defparam add_1176_5.INIT1 = 16'hf555;
    defparam add_1176_5.INJECT1_0 = "NO";
    defparam add_1176_5.INJECT1_1 = "NO";
    LUT4 i18266_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut_4_lut (.A(n21893), .B(ss[0]), 
         .C(ss[2]), .D(ss[1]), .Z(n20582)) /* synthesis lut_function=(!(A+(B (C (D))+!B !(C+(D))))) */ ;
    defparam i18266_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut_4_lut.init = 16'h1554;
    CCU2D add_191_11 (.A0(Out3[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18710), 
          .COUT(n18711), .S0(n1208[9]), .S1(n1208[10]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_11.INIT0 = 16'h5aaa;
    defparam add_191_11.INIT1 = 16'h5aaa;
    defparam add_191_11.INJECT1_0 = "NO";
    defparam add_191_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_457_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(ss[3]), 
         .D(n22388), .Z(n21877)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_457_3_lut_4_lut.init = 16'h0006;
    PFUMX mux_1802_i1 (.BLUT(subIn2_24__N_1301[0]), .ALUT(subIn2_24__N_1114[0]), 
          .C0(n20586), .Z(subIn2[0]));
    LUT4 i1815_1_lut_rep_477 (.A(ss[0]), .Z(n21897)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1815_1_lut_rep_477.init = 16'h5555;
    LUT4 i1_2_lut_4_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(n21922), .D(n22388), 
         .Z(n4148)) /* synthesis lut_function=(!(A+(B (C+(D))+!B ((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h0014;
    CCU2D add_1180_9 (.A0(n5152), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5154), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18674), 
          .COUT(n18675), .S0(n2245[7]), .S1(n2245[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_9.INIT0 = 16'hf555;
    defparam add_1180_9.INIT1 = 16'hf555;
    defparam add_1180_9.INJECT1_0 = "NO";
    defparam add_1180_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_478 (.A(ss[0]), .B(ss[3]), .Z(n21898)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_rep_478.init = 16'h8888;
    CCU2D add_1180_7 (.A0(n5148), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5150), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18673), 
          .COUT(n18674), .S0(n2245[5]), .S1(n2245[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_7.INIT0 = 16'hf555;
    defparam add_1180_7.INIT1 = 16'hf555;
    defparam add_1180_7.INJECT1_0 = "NO";
    defparam add_1180_7.INJECT1_1 = "NO";
    LUT4 i7_4_lut_adj_120 (.A(Out2[3]), .B(n14_adj_1862), .C(n10_adj_1863), 
         .D(Out2[4]), .Z(n19127)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam i7_4_lut_adj_120.init = 16'hfffe;
    LUT4 i6_4_lut_adj_121 (.A(Out2[11]), .B(Out2[7]), .C(Out2[2]), .D(Out2[10]), 
         .Z(n14_adj_1862)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam i6_4_lut_adj_121.init = 16'hfffe;
    LUT4 i2_2_lut_adj_122 (.A(Out2[9]), .B(Out2[1]), .Z(n10_adj_1863)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam i2_2_lut_adj_122.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n20055)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(204[2] 392[9])
    defparam i1_2_lut_3_lut.init = 16'h0808;
    PFUMX mux_140_i25 (.BLUT(n558[24]), .ALUT(n678[24]), .C0(n20525), 
          .Z(addIn2_28__N_1337[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i17 (.BLUT(n558[16]), .ALUT(n678[16]), .C0(n20525), 
          .Z(addIn2_28__N_1337[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i7 (.BLUT(n558[6]), .ALUT(n678[6]), .C0(n20525), .Z(addIn2_28__N_1337[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i4_4_lut_adj_123 (.A(Out2[5]), .B(Out2[6]), .C(Out2[0]), .D(n6_adj_1864), 
         .Z(n19128)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam i4_4_lut_adj_123.init = 16'hfffe;
    LUT4 i1_2_lut_adj_124 (.A(Out2[8]), .B(Out2[12]), .Z(n6_adj_1864)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam i1_2_lut_adj_124.init = 16'heeee;
    PFUMX mux_140_i26 (.BLUT(n558[25]), .ALUT(n678[25]), .C0(n20525), 
          .Z(addIn2_28__N_1337[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i18 (.BLUT(n558[17]), .ALUT(n678[17]), .C0(n20525), 
          .Z(addIn2_28__N_1337[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1_2_lut_rep_483 (.A(ss[0]), .B(ss[3]), .Z(n21903)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_483.init = 16'hbbbb;
    PFUMX mux_140_i8 (.BLUT(n558[7]), .ALUT(n678[7]), .C0(n20525), .Z(addIn2_28__N_1337[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1_2_lut_3_lut_adj_125 (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n20202)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_3_lut_adj_125.init = 16'hfbfb;
    CCU2D add_1176_3 (.A0(n1187[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18771), 
          .COUT(n18772), .S0(n2177[1]), .S1(n2177[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(343[20:29])
    defparam add_1176_3.INIT0 = 16'hf555;
    defparam add_1176_3.INIT1 = 16'hf555;
    defparam add_1176_3.INJECT1_0 = "NO";
    defparam add_1176_3.INJECT1_1 = "NO";
    CCU2D add_191_9 (.A0(Out3[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18709), 
          .COUT(n18710), .S0(n1208[7]), .S1(n1208[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_9.INIT0 = 16'h5aaa;
    defparam add_191_9.INIT1 = 16'h5aaa;
    defparam add_191_9.INJECT1_0 = "NO";
    defparam add_191_9.INJECT1_1 = "NO";
    CCU2D add_191_7 (.A0(Out3[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18708), 
          .COUT(n18709), .S0(n1208[5]), .S1(n1208[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_7.INIT0 = 16'h5aaa;
    defparam add_191_7.INIT1 = 16'h5aaa;
    defparam add_191_7.INJECT1_0 = "NO";
    defparam add_191_7.INJECT1_1 = "NO";
    PFUMX mux_140_i27 (.BLUT(n558[26]), .ALUT(n678[26]), .C0(n20525), 
          .Z(addIn2_28__N_1337[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1176_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18771), 
          .S1(n2177[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(343[20:29])
    defparam add_1176_1.INIT0 = 16'hF000;
    defparam add_1176_1.INIT1 = 16'h0aaa;
    defparam add_1176_1.INJECT1_0 = "NO";
    defparam add_1176_1.INJECT1_1 = "NO";
    CCU2D add_191_5 (.A0(Out3[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18707), 
          .COUT(n18708), .S0(n1208[3]), .S1(n1208[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_5.INIT0 = 16'h5aaa;
    defparam add_191_5.INIT1 = 16'h5aaa;
    defparam add_191_5.INJECT1_0 = "NO";
    defparam add_191_5.INJECT1_1 = "NO";
    CCU2D add_191_3 (.A0(Out3[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18706), 
          .COUT(n18707), .S0(n1208[1]), .S1(n1208[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_3.INIT0 = 16'h5aaa;
    defparam add_191_3.INIT1 = 16'h5aaa;
    defparam add_191_3.INJECT1_0 = "NO";
    defparam add_191_3.INJECT1_1 = "NO";
    PFUMX mux_140_i19 (.BLUT(n558[18]), .ALUT(n678[18]), .C0(n20525), 
          .Z(addIn2_28__N_1337[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i9 (.BLUT(n558[8]), .ALUT(n678[8]), .C0(n20525), .Z(addIn2_28__N_1337[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i28 (.BLUT(n558[27]), .ALUT(n678[27]), .C0(n20525), 
          .Z(addIn2_28__N_1337[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D addOut_2064_add_4_29 (.A0(multOut[27]), .B0(n16286), .C0(addOut[27]), 
          .D0(addIn2_28__N_1207[27]), .A1(multOut[28]), .B1(n16286), .C1(addOut[28]), 
          .D1(addIn2_28__N_1207[28]), .CIN(n18834), .S0(n121[27]), .S1(n121[28]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_29.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_29.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_29.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_29.INJECT1_1 = "NO";
    PFUMX mux_140_i20 (.BLUT(n558[19]), .ALUT(n678[19]), .C0(n20525), 
          .Z(addIn2_28__N_1337[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1175_11 (.A0(n1166[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18770), 
          .S0(n2165[9]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(335[20:29])
    defparam add_1175_11.INIT0 = 16'hf555;
    defparam add_1175_11.INIT1 = 16'h0000;
    defparam add_1175_11.INJECT1_0 = "NO";
    defparam add_1175_11.INJECT1_1 = "NO";
    CCU2D add_191_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[13]), .B1(n19124), .C1(n19125), .D1(Out3[28]), .COUT(n18706), 
          .S1(n1208[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(317[17:21])
    defparam add_191_1.INIT0 = 16'hF000;
    defparam add_191_1.INIT1 = 16'h56aa;
    defparam add_191_1.INJECT1_0 = "NO";
    defparam add_191_1.INJECT1_1 = "NO";
    CCU2D add_1180_5 (.A0(n5144), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5146), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18672), 
          .COUT(n18673), .S0(n2245[3]), .S1(n2245[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_5.INIT0 = 16'hf555;
    defparam add_1180_5.INIT1 = 16'hf555;
    defparam add_1180_5.INJECT1_0 = "NO";
    defparam add_1180_5.INJECT1_1 = "NO";
    PFUMX mux_140_i10 (.BLUT(n558[9]), .ALUT(n678[9]), .C0(n20525), .Z(addIn2_28__N_1337[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1180_3 (.A0(n5140), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5142), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18671), 
          .COUT(n18672), .S0(n2245[1]), .S1(n2245[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(126[13] 142[6])
    defparam add_1180_3.INIT0 = 16'hf555;
    defparam add_1180_3.INIT1 = 16'hf555;
    defparam add_1180_3.INJECT1_0 = "NO";
    defparam add_1180_3.INJECT1_1 = "NO";
    PFUMX mux_140_i11 (.BLUT(n558[10]), .ALUT(n678[10]), .C0(n20525), 
          .Z(addIn2_28__N_1337[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D addOut_2064_add_4_27 (.A0(multOut[25]), .B0(n16286), .C0(addOut[25]), 
          .D0(addIn2_28__N_1207[25]), .A1(multOut[26]), .B1(n16286), .C1(addOut[26]), 
          .D1(addIn2_28__N_1207[26]), .CIN(n18833), .COUT(n18834), .S0(n121[25]), 
          .S1(n121[26]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_27.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_27.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_27.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_27.INJECT1_1 = "NO";
    CCU2D add_187_17 (.A0(Out2[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18705), 
          .S0(n1187[15]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_17.INIT0 = 16'h5aaa;
    defparam add_187_17.INIT1 = 16'h0000;
    defparam add_187_17.INJECT1_0 = "NO";
    defparam add_187_17.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_25 (.A0(multOut[23]), .B0(n16286), .C0(addOut[23]), 
          .D0(addIn2_28__N_1207[23]), .A1(multOut[24]), .B1(n16286), .C1(addOut[24]), 
          .D1(addIn2_28__N_1207[24]), .CIN(n18832), .COUT(n18833), .S0(n121[23]), 
          .S1(n121[24]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_25.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_25.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_25.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_25.INJECT1_1 = "NO";
    CCU2D add_16119_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18920), 
          .S0(n920));
    defparam add_16119_cout.INIT0 = 16'h0000;
    defparam add_16119_cout.INIT1 = 16'h0000;
    defparam add_16119_cout.INJECT1_0 = "NO";
    defparam add_16119_cout.INJECT1_1 = "NO";
    PFUMX mux_140_i29 (.BLUT(n558[28]), .ALUT(n678[28]), .C0(n20525), 
          .Z(addIn2_28__N_1337[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_16119_22 (.A0(addOut[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18919), .COUT(n18920));
    defparam add_16119_22.INIT0 = 16'h5555;
    defparam add_16119_22.INIT1 = 16'hf555;
    defparam add_16119_22.INJECT1_0 = "NO";
    defparam add_16119_22.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_23 (.A0(multOut[21]), .B0(n16286), .C0(addOut[21]), 
          .D0(addIn2_28__N_1207[21]), .A1(multOut[22]), .B1(n16286), .C1(addOut[22]), 
          .D1(addIn2_28__N_1207[22]), .CIN(n18831), .COUT(n18832), .S0(n121[21]), 
          .S1(n121[22]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_23.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_23.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_23.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_23.INJECT1_1 = "NO";
    CCU2D add_1175_9 (.A0(n1166[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18769), 
          .COUT(n18770), .S0(n2165[7]), .S1(n2165[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(335[20:29])
    defparam add_1175_9.INIT0 = 16'hf555;
    defparam add_1175_9.INIT1 = 16'hf555;
    defparam add_1175_9.INJECT1_0 = "NO";
    defparam add_1175_9.INJECT1_1 = "NO";
    CCU2D add_187_15 (.A0(Out2[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18704), 
          .COUT(n18705), .S0(n1187[13]), .S1(n1187[14]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_15.INIT0 = 16'h5aaa;
    defparam add_187_15.INIT1 = 16'h5aaa;
    defparam add_187_15.INJECT1_0 = "NO";
    defparam add_187_15.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_21 (.A0(multOut[19]), .B0(n16286), .C0(addOut[19]), 
          .D0(addIn2_28__N_1207[19]), .A1(multOut[20]), .B1(n16286), .C1(addOut[20]), 
          .D1(addIn2_28__N_1207[20]), .CIN(n18830), .COUT(n18831), .S0(n121[19]), 
          .S1(n121[20]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_21.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_21.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_21.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_21.INJECT1_1 = "NO";
    CCU2D add_16119_20 (.A0(addOut[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18918), .COUT(n18919));
    defparam add_16119_20.INIT0 = 16'h5555;
    defparam add_16119_20.INIT1 = 16'h5555;
    defparam add_16119_20.INJECT1_0 = "NO";
    defparam add_16119_20.INJECT1_1 = "NO";
    CCU2D add_187_13 (.A0(Out2[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18703), 
          .COUT(n18704), .S0(n1187[11]), .S1(n1187[12]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_13.INIT0 = 16'h5aaa;
    defparam add_187_13.INIT1 = 16'h5aaa;
    defparam add_187_13.INJECT1_0 = "NO";
    defparam add_187_13.INJECT1_1 = "NO";
    LUT4 i1755_1_lut (.A(n42), .Z(subIn1_24__N_1300)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(137[34:50])
    defparam i1755_1_lut.init = 16'h5555;
    CCU2D addOut_2064_add_4_19 (.A0(multOut[17]), .B0(n16286), .C0(addOut[17]), 
          .D0(addIn2_28__N_1207[17]), .A1(multOut[18]), .B1(n16286), .C1(addOut[18]), 
          .D1(addIn2_28__N_1207[18]), .CIN(n18829), .COUT(n18830), .S0(n121[17]), 
          .S1(n121[18]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_19.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_19.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_19.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_19.INJECT1_1 = "NO";
    PFUMX mux_140_i21 (.BLUT(n558[20]), .ALUT(n678[20]), .C0(n20525), 
          .Z(addIn2_28__N_1337[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i12 (.BLUT(n558[11]), .ALUT(n678[11]), .C0(n20525), 
          .Z(addIn2_28__N_1337[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i22 (.BLUT(n558[21]), .ALUT(n678[21]), .C0(n20525), 
          .Z(addIn2_28__N_1337[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i13560_3_lut_4_lut (.A(n920), .B(n3636), .C(n22388), .D(addOut[6]), 
         .Z(intgOut0_28__N_735[6])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i13560_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i1756_1_lut (.A(n49), .Z(dirout_m3_N_1578)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(139[35:51])
    defparam i1756_1_lut.init = 16'h5555;
    PFUMX mux_140_i13 (.BLUT(n558[12]), .ALUT(n678[12]), .C0(n20525), 
          .Z(addIn2_28__N_1337[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1754_1_lut (.A(n35), .Z(subIn1_24__N_1113)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(135[34:50])
    defparam i1754_1_lut.init = 16'h5555;
    PFUMX mux_140_i14 (.BLUT(n558[13]), .ALUT(n678[13]), .C0(n20525), 
          .Z(addIn2_28__N_1337[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i23 (.BLUT(n558[22]), .ALUT(n678[22]), .C0(n20525), 
          .Z(addIn2_28__N_1337[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i24 (.BLUT(n558[23]), .ALUT(n678[23]), .C0(n20525), 
          .Z(addIn2_28__N_1337[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_140_i15 (.BLUT(n558[14]), .ALUT(n678[14]), .C0(n20525), 
          .Z(addIn2_28__N_1337[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1757_1_lut (.A(n56), .Z(dirout_m4_N_1581)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(141[35:51])
    defparam i1757_1_lut.init = 16'h5555;
    PFUMX mux_140_i16 (.BLUT(n558[15]), .ALUT(n678[15]), .C0(n20525), 
          .Z(addIn2_28__N_1337[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D addOut_2064_add_4_17 (.A0(multOut[15]), .B0(n16286), .C0(addOut[15]), 
          .D0(addIn2_28__N_1207[15]), .A1(multOut[16]), .B1(n16286), .C1(addOut[16]), 
          .D1(addIn2_28__N_1207[16]), .CIN(n18828), .COUT(n18829), .S0(n121[15]), 
          .S1(n121[16]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_17.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_17.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_17.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_17.INJECT1_1 = "NO";
    CCU2D add_1175_7 (.A0(n1166[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18768), 
          .COUT(n18769), .S0(n2165[5]), .S1(n2165[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(335[20:29])
    defparam add_1175_7.INIT0 = 16'hf555;
    defparam add_1175_7.INIT1 = 16'hf555;
    defparam add_1175_7.INJECT1_0 = "NO";
    defparam add_1175_7.INJECT1_1 = "NO";
    CCU2D add_187_11 (.A0(Out2[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18702), 
          .COUT(n18703), .S0(n1187[9]), .S1(n1187[10]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_11.INIT0 = 16'h5aaa;
    defparam add_187_11.INIT1 = 16'h5aaa;
    defparam add_187_11.INJECT1_0 = "NO";
    defparam add_187_11.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_15 (.A0(multOut[13]), .B0(n16286), .C0(addOut[13]), 
          .D0(addIn2_28__N_1207[13]), .A1(multOut[14]), .B1(n16286), .C1(addOut[14]), 
          .D1(addIn2_28__N_1207[14]), .CIN(n18827), .COUT(n18828), .S0(n121[13]), 
          .S1(n121[14]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_15.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_15.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_15.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_15.INJECT1_1 = "NO";
    CCU2D add_16119_18 (.A0(addOut[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18917), .COUT(n18918));
    defparam add_16119_18.INIT0 = 16'h5555;
    defparam add_16119_18.INIT1 = 16'h5555;
    defparam add_16119_18.INJECT1_0 = "NO";
    defparam add_16119_18.INJECT1_1 = "NO";
    CCU2D add_1175_5 (.A0(n1166[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18767), 
          .COUT(n18768), .S0(n2165[3]), .S1(n2165[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(335[20:29])
    defparam add_1175_5.INIT0 = 16'hf555;
    defparam add_1175_5.INIT1 = 16'hf555;
    defparam add_1175_5.INJECT1_0 = "NO";
    defparam add_1175_5.INJECT1_1 = "NO";
    CCU2D add_187_9 (.A0(Out2[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18701), 
          .COUT(n18702), .S0(n1187[7]), .S1(n1187[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_9.INIT0 = 16'h5aaa;
    defparam add_187_9.INIT1 = 16'h5aaa;
    defparam add_187_9.INJECT1_0 = "NO";
    defparam add_187_9.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_13 (.A0(multOut[11]), .B0(n16286), .C0(addOut[11]), 
          .D0(addIn2_28__N_1207[11]), .A1(multOut[12]), .B1(n16286), .C1(addOut[12]), 
          .D1(addIn2_28__N_1207[12]), .CIN(n18826), .COUT(n18827), .S0(n121[11]), 
          .S1(n121[12]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_13.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_13.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_13.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_13.INJECT1_1 = "NO";
    CCU2D add_16119_16 (.A0(addOut[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18916), .COUT(n18917));
    defparam add_16119_16.INIT0 = 16'h5555;
    defparam add_16119_16.INIT1 = 16'h5555;
    defparam add_16119_16.INJECT1_0 = "NO";
    defparam add_16119_16.INJECT1_1 = "NO";
    CCU2D add_187_7 (.A0(Out2[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18700), 
          .COUT(n18701), .S0(n1187[5]), .S1(n1187[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_7.INIT0 = 16'h5aaa;
    defparam add_187_7.INIT1 = 16'h5aaa;
    defparam add_187_7.INJECT1_0 = "NO";
    defparam add_187_7.INJECT1_1 = "NO";
    CCU2D add_1175_3 (.A0(n1166[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18766), 
          .COUT(n18767), .S0(n2165[1]), .S1(n2165[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(335[20:29])
    defparam add_1175_3.INIT0 = 16'hf555;
    defparam add_1175_3.INIT1 = 16'hf555;
    defparam add_1175_3.INJECT1_0 = "NO";
    defparam add_1175_3.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_11 (.A0(multOut[9]), .B0(n16286), .C0(addOut[9]), 
          .D0(addIn2_28__N_1207[9]), .A1(multOut[10]), .B1(n16286), .C1(addOut[10]), 
          .D1(addIn2_28__N_1207[10]), .CIN(n18825), .COUT(n18826), .S0(n121[9]), 
          .S1(n121[10]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_11.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_11.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_11.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_11.INJECT1_1 = "NO";
    CCU2D add_1175_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18766), 
          .S1(n2165[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(335[20:29])
    defparam add_1175_1.INIT0 = 16'hF000;
    defparam add_1175_1.INIT1 = 16'h0aaa;
    defparam add_1175_1.INJECT1_0 = "NO";
    defparam add_1175_1.INJECT1_1 = "NO";
    LUT4 mux_205_i4_3_lut_4_lut_3_lut (.A(n30_c), .B(n1166[15]), .C(n2165[3]), 
         .Z(n1302[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(334[25:42])
    defparam mux_205_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    PFUMX mux_137_i24 (.BLUT(n588[23]), .ALUT(intgOut3_c[23]), .C0(n21835), 
          .Z(n618[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i25 (.BLUT(n588[24]), .ALUT(intgOut3_c[24]), .C0(n21835), 
          .Z(n618[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i26 (.BLUT(n588[25]), .ALUT(intgOut3_c[25]), .C0(n21835), 
          .Z(n618[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i27 (.BLUT(n588[26]), .ALUT(intgOut3_c[26]), .C0(n21835), 
          .Z(n618[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i28 (.BLUT(n588[27]), .ALUT(intgOut3_c[27]), .C0(n21835), 
          .Z(n618[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_187_5 (.A0(Out2[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18699), 
          .COUT(n18700), .S0(n1187[3]), .S1(n1187[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_5.INIT0 = 16'h5aaa;
    defparam add_187_5.INIT1 = 16'h5aaa;
    defparam add_187_5.INJECT1_0 = "NO";
    defparam add_187_5.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_9 (.A0(multOut[7]), .B0(n16286), .C0(addOut[7]), 
          .D0(addIn2_28__N_1207[7]), .A1(multOut[8]), .B1(n16286), .C1(addOut[8]), 
          .D1(addIn2_28__N_1207[8]), .CIN(n18824), .COUT(n18825), .S0(n121[7]), 
          .S1(n121[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_9.INIT0 = 16'h569a;
    defparam addOut_2064_add_4_9.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_9.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_9.INJECT1_1 = "NO";
    PFUMX mux_137_i7 (.BLUT(n588[6]), .ALUT(intgOut3_c[6]), .C0(n21835), 
          .Z(n618[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_16119_14 (.A0(addOut[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18915), .COUT(n18916));
    defparam add_16119_14.INIT0 = 16'h5aaa;
    defparam add_16119_14.INIT1 = 16'h5555;
    defparam add_16119_14.INJECT1_0 = "NO";
    defparam add_16119_14.INJECT1_1 = "NO";
    PFUMX mux_137_i29 (.BLUT(n588[28]), .ALUT(intgOut3_c[28]), .C0(n21835), 
          .Z(n618[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i8 (.BLUT(n588[7]), .ALUT(intgOut3_c[7]), .C0(n21835), 
          .Z(n618[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i9 (.BLUT(n588[8]), .ALUT(intgOut3_c[8]), .C0(n21835), 
          .Z(n618[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1_2_lut_rep_399_4_lut_4_lut (.A(n21835), .B(n35), .C(n21867), 
         .D(n21866), .Z(n21819)) /* synthesis lut_function=(A (B)+!A !((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(171[9:16])
    defparam i1_2_lut_rep_399_4_lut_4_lut.init = 16'h888c;
    PFUMX mux_137_i10 (.BLUT(n588[9]), .ALUT(intgOut3_c[9]), .C0(n21835), 
          .Z(n618[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i11 (.BLUT(n588[10]), .ALUT(intgOut3_c[10]), .C0(n21835), 
          .Z(n618[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i12 (.BLUT(n588[11]), .ALUT(intgOut3_c[11]), .C0(n21835), 
          .Z(n618[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i13 (.BLUT(n588[12]), .ALUT(intgOut3_c[12]), .C0(n21835), 
          .Z(n618[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i14 (.BLUT(n588[13]), .ALUT(intgOut3_c[13]), .C0(n21835), 
          .Z(n618[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D sub_17_rep_2_add_2_23 (.A0(n2245[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18764), .S0(n4183), .S1(n4182));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_23.INIT0 = 16'h5555;
    defparam sub_17_rep_2_add_2_23.INIT1 = 16'h5555;
    defparam sub_17_rep_2_add_2_23.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_23.INJECT1_1 = "NO";
    CCU2D add_187_3 (.A0(Out2[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18698), 
          .COUT(n18699), .S0(n1187[1]), .S1(n1187[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_3.INIT0 = 16'h5aaa;
    defparam add_187_3.INIT1 = 16'h5aaa;
    defparam add_187_3.INJECT1_0 = "NO";
    defparam add_187_3.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_7 (.A0(multOut[5]), .B0(n16286), .C0(n13), 
          .D0(addOut[5]), .A1(multOut[6]), .B1(n16286), .C1(addOut[6]), 
          .D1(addIn2_28__N_1207[6]), .CIN(n18823), .COUT(n18824), .S0(n121[5]), 
          .S1(n121[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_7.INIT0 = 16'h596a;
    defparam addOut_2064_add_4_7.INIT1 = 16'h569a;
    defparam addOut_2064_add_4_7.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_7.INJECT1_1 = "NO";
    CCU2D add_16119_12 (.A0(addOut[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18914), .COUT(n18915));
    defparam add_16119_12.INIT0 = 16'h5aaa;
    defparam add_16119_12.INIT1 = 16'h5aaa;
    defparam add_16119_12.INJECT1_0 = "NO";
    defparam add_16119_12.INJECT1_1 = "NO";
    CCU2D add_187_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[13]), .B1(n19127), .C1(n19128), .D1(Out2[28]), .COUT(n18698), 
          .S1(n1187[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(316[17:21])
    defparam add_187_1.INIT0 = 16'hF000;
    defparam add_187_1.INIT1 = 16'h56aa;
    defparam add_187_1.INJECT1_0 = "NO";
    defparam add_187_1.INJECT1_1 = "NO";
    CCU2D sub_17_rep_2_add_2_21 (.A0(n2245[19]), .B0(n7), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18763), .COUT(n18764), .S0(n4185), .S1(n4184));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_21.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_21.INIT1 = 16'h5555;
    defparam sub_17_rep_2_add_2_21.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_21.INJECT1_1 = "NO";
    PFUMX mux_137_i15 (.BLUT(n588[14]), .ALUT(intgOut3_c[14]), .C0(n21835), 
          .Z(n618[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D addOut_2064_add_4_5 (.A0(multOut[3]), .B0(n16286), .C0(n13_adj_9), 
          .D0(addOut[3]), .A1(multOut[4]), .B1(n16286), .C1(n13_adj_10), 
          .D1(addOut[4]), .CIN(n18822), .COUT(n18823), .S0(n121[3]), 
          .S1(n121[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_5.INIT0 = 16'h596a;
    defparam addOut_2064_add_4_5.INIT1 = 16'h596a;
    defparam addOut_2064_add_4_5.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_5.INJECT1_1 = "NO";
    CCU2D sub_17_rep_2_add_2_19 (.A0(n2245[17]), .B0(subIn2[17]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[18]), .B1(subIn2[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18762), .COUT(n18763), .S0(n4187), .S1(n4186));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_19.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_19.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_19.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_19.INJECT1_1 = "NO";
    CCU2D add_183_17 (.A0(Out1[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18697), 
          .S0(n1166[15]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_17.INIT0 = 16'h5aaa;
    defparam add_183_17.INIT1 = 16'h0000;
    defparam add_183_17.INJECT1_0 = "NO";
    defparam add_183_17.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_3 (.A0(multOut[1]), .B0(n16286), .C0(n13_adj_11), 
          .D0(addOut[1]), .A1(multOut[2]), .B1(n16286), .C1(n13_adj_12), 
          .D1(addOut[2]), .CIN(n18821), .COUT(n18822), .S0(n121[1]), 
          .S1(n121[2]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_3.INIT0 = 16'h596a;
    defparam addOut_2064_add_4_3.INIT1 = 16'h596a;
    defparam addOut_2064_add_4_3.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_3.INJECT1_1 = "NO";
    CCU2D add_16119_10 (.A0(addOut[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18913), .COUT(n18914));
    defparam add_16119_10.INIT0 = 16'h5555;
    defparam add_16119_10.INIT1 = 16'h5aaa;
    defparam add_16119_10.INJECT1_0 = "NO";
    defparam add_16119_10.INJECT1_1 = "NO";
    CCU2D sub_17_rep_2_add_2_17 (.A0(n2245[15]), .B0(subIn2[15]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[16]), .B1(subIn2[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18761), .COUT(n18762), .S0(n4189), .S1(n4188));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_17.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_17.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_17.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_17.INJECT1_1 = "NO";
    CCU2D add_183_15 (.A0(Out1[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18696), 
          .COUT(n18697), .S0(n1166[13]), .S1(n1166[14]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_15.INIT0 = 16'h5aaa;
    defparam add_183_15.INIT1 = 16'h5aaa;
    defparam add_183_15.INJECT1_0 = "NO";
    defparam add_183_15.INJECT1_1 = "NO";
    CCU2D addOut_2064_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(multOut[0]), .B1(n16286), .C1(n14), .D1(addOut[0]), 
          .COUT(n18821), .S1(n121[0]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064_add_4_1.INIT0 = 16'hF000;
    defparam addOut_2064_add_4_1.INIT1 = 16'h596a;
    defparam addOut_2064_add_4_1.INJECT1_0 = "NO";
    defparam addOut_2064_add_4_1.INJECT1_1 = "NO";
    CCU2D add_16119_8 (.A0(addOut[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18912), .COUT(n18913));
    defparam add_16119_8.INIT0 = 16'h5555;
    defparam add_16119_8.INIT1 = 16'h5aaa;
    defparam add_16119_8.INJECT1_0 = "NO";
    defparam add_16119_8.INJECT1_1 = "NO";
    CCU2D add_183_13 (.A0(Out1[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18695), 
          .COUT(n18696), .S0(n1166[11]), .S1(n1166[12]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_13.INIT0 = 16'h5aaa;
    defparam add_183_13.INIT1 = 16'h5aaa;
    defparam add_183_13.INJECT1_0 = "NO";
    defparam add_183_13.INJECT1_1 = "NO";
    PFUMX mux_137_i16 (.BLUT(n588[15]), .ALUT(intgOut3_c[15]), .C0(n21835), 
          .Z(n618[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1_2_lut_rep_502 (.A(n22379), .B(ss[1]), .Z(n21922)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_502.init = 16'heeee;
    LUT4 i1_3_lut_rep_450_4_lut (.A(ss[2]), .B(ss[1]), .C(ss[3]), .D(n22388), 
         .Z(n21870)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i1_3_lut_rep_450_4_lut.init = 16'h001e;
    PFUMX mux_137_i17 (.BLUT(n588[16]), .ALUT(intgOut3_c[16]), .C0(n21835), 
          .Z(n618[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D sub_17_rep_2_add_2_15 (.A0(n2245[13]), .B0(subIn2[13]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[14]), .B1(subIn2[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18760), .COUT(n18761), .S0(n4191), .S1(n4190));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_15.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_15.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_15.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_503 (.A(ss[0]), .B(ss[3]), .Z(n21923)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_503.init = 16'heeee;
    FD1S3AX addOut_2064__i1 (.D(n121[1]), .CK(clk_N_683), .Q(addOut[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i1.GSR = "ENABLED";
    LUT4 i2_2_lut_rep_465_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), 
         .D(n22379), .Z(n21885)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(235[3] 390[12])
    defparam i2_2_lut_rep_465_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_504 (.A(ss[0]), .B(ss[2]), .Z(n21924)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_504.init = 16'h8888;
    CCU2D sub_17_rep_2_add_2_13 (.A0(n2245[11]), .B0(subIn2[11]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[12]), .B1(subIn2[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18759), .COUT(n18760), .S0(n4193), .S1(n4192));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_13.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_13.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_13.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_13.INJECT1_1 = "NO";
    PFUMX mux_137_i18 (.BLUT(n588[17]), .ALUT(intgOut3_c[17]), .C0(n21835), 
          .Z(n618[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i19 (.BLUT(n588[18]), .ALUT(intgOut3_c[18]), .C0(n21835), 
          .Z(n618[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX i18454 (.BLUT(n21931), .ALUT(n21932), .C0(ss[2]), .Z(n21933));
    PFUMX mux_137_i20 (.BLUT(n588[19]), .ALUT(intgOut3_c[19]), .C0(n21835), 
          .Z(n618[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i21 (.BLUT(n588[20]), .ALUT(intgOut3_c[20]), .C0(n21835), 
          .Z(n618[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX mux_137_i22 (.BLUT(n588[21]), .ALUT(intgOut3_c[21]), .C0(n21835), 
          .Z(n618[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    PFUMX i18452 (.BLUT(n21928), .ALUT(n21929), .C0(ss[0]), .Z(n4133));
    PFUMX mux_137_i23 (.BLUT(n588[22]), .ALUT(intgOut3_c[22]), .C0(n21835), 
          .Z(n618[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    FD1S3AX addOut_2064__i2 (.D(n121[2]), .CK(clk_N_683), .Q(addOut[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i2.GSR = "ENABLED";
    FD1S3AX addOut_2064__i3 (.D(n121[3]), .CK(clk_N_683), .Q(addOut[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i3.GSR = "ENABLED";
    FD1S3AX addOut_2064__i4 (.D(n121[4]), .CK(clk_N_683), .Q(addOut[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i4.GSR = "ENABLED";
    FD1S3AX addOut_2064__i5 (.D(n121[5]), .CK(clk_N_683), .Q(addOut[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i5.GSR = "ENABLED";
    FD1S3AX addOut_2064__i6 (.D(n121[6]), .CK(clk_N_683), .Q(addOut[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i6.GSR = "ENABLED";
    FD1S3AX addOut_2064__i7 (.D(n121[7]), .CK(clk_N_683), .Q(addOut[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i7.GSR = "ENABLED";
    FD1S3AX addOut_2064__i8 (.D(n121[8]), .CK(clk_N_683), .Q(addOut[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i8.GSR = "ENABLED";
    FD1S3AX addOut_2064__i9 (.D(n121[9]), .CK(clk_N_683), .Q(addOut[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i9.GSR = "ENABLED";
    FD1S3AX addOut_2064__i10 (.D(n121[10]), .CK(clk_N_683), .Q(addOut[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i10.GSR = "ENABLED";
    FD1S3AX addOut_2064__i11 (.D(n121[11]), .CK(clk_N_683), .Q(addOut[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i11.GSR = "ENABLED";
    FD1S3AX addOut_2064__i12 (.D(n121[12]), .CK(clk_N_683), .Q(addOut[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i12.GSR = "ENABLED";
    FD1S3AX addOut_2064__i13 (.D(n121[13]), .CK(clk_N_683), .Q(addOut[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i13.GSR = "ENABLED";
    FD1S3AX addOut_2064__i14 (.D(n121[14]), .CK(clk_N_683), .Q(addOut[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i14.GSR = "ENABLED";
    FD1S3AX addOut_2064__i15 (.D(n121[15]), .CK(clk_N_683), .Q(addOut[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i15.GSR = "ENABLED";
    FD1S3AX addOut_2064__i16 (.D(n121[16]), .CK(clk_N_683), .Q(addOut[16])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i16.GSR = "ENABLED";
    FD1S3AX addOut_2064__i17 (.D(n121[17]), .CK(clk_N_683), .Q(addOut[17])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i17.GSR = "ENABLED";
    FD1S3AX addOut_2064__i18 (.D(n121[18]), .CK(clk_N_683), .Q(addOut[18])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i18.GSR = "ENABLED";
    FD1S3AX addOut_2064__i19 (.D(n121[19]), .CK(clk_N_683), .Q(addOut[19])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i19.GSR = "ENABLED";
    FD1S3AX addOut_2064__i20 (.D(n121[20]), .CK(clk_N_683), .Q(addOut[20])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i20.GSR = "ENABLED";
    FD1S3AX addOut_2064__i21 (.D(n121[21]), .CK(clk_N_683), .Q(addOut[21])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i21.GSR = "ENABLED";
    FD1S3AX addOut_2064__i22 (.D(n121[22]), .CK(clk_N_683), .Q(addOut[22])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i22.GSR = "ENABLED";
    FD1S3AX addOut_2064__i23 (.D(n121[23]), .CK(clk_N_683), .Q(addOut[23])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i23.GSR = "ENABLED";
    FD1S3AX addOut_2064__i24 (.D(n121[24]), .CK(clk_N_683), .Q(addOut[24])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i24.GSR = "ENABLED";
    FD1S3AX addOut_2064__i25 (.D(n121[25]), .CK(clk_N_683), .Q(addOut[25])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i25.GSR = "ENABLED";
    FD1S3AX addOut_2064__i26 (.D(n121[26]), .CK(clk_N_683), .Q(addOut[26])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i26.GSR = "ENABLED";
    FD1S3AX addOut_2064__i27 (.D(n121[27]), .CK(clk_N_683), .Q(addOut[27])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i27.GSR = "ENABLED";
    FD1S3AX addOut_2064__i28 (.D(n121[28]), .CK(clk_N_683), .Q(addOut[28])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(230[13:19])
    defparam addOut_2064__i28.GSR = "ENABLED";
    CCU2D add_183_11 (.A0(Out1[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18694), 
          .COUT(n18695), .S0(n1166[9]), .S1(n1166[10]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_11.INIT0 = 16'h5aaa;
    defparam add_183_11.INIT1 = 16'h5aaa;
    defparam add_183_11.INJECT1_0 = "NO";
    defparam add_183_11.INJECT1_1 = "NO";
    CCU2D add_16119_6 (.A0(addOut[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18911), .COUT(n18912));
    defparam add_16119_6.INIT0 = 16'h5555;
    defparam add_16119_6.INIT1 = 16'h5555;
    defparam add_16119_6.INJECT1_0 = "NO";
    defparam add_16119_6.INJECT1_1 = "NO";
    CCU2D sub_17_rep_2_add_2_11 (.A0(n2245[9]), .B0(subIn2[9]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[10]), .B1(subIn2[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18758), .COUT(n18759), .S0(n4195), .S1(n4194));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_11.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_11.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_11.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_11.INJECT1_1 = "NO";
    CCU2D add_183_9 (.A0(Out1[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18693), 
          .COUT(n18694), .S0(n1166[7]), .S1(n1166[8]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_9.INIT0 = 16'h5aaa;
    defparam add_183_9.INIT1 = 16'h5aaa;
    defparam add_183_9.INJECT1_0 = "NO";
    defparam add_183_9.INJECT1_1 = "NO";
    CCU2D add_16119_4 (.A0(addOut[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18910), .COUT(n18911));
    defparam add_16119_4.INIT0 = 16'h5aaa;
    defparam add_16119_4.INIT1 = 16'h5555;
    defparam add_16119_4.INJECT1_0 = "NO";
    defparam add_16119_4.INJECT1_1 = "NO";
    CCU2D add_183_7 (.A0(Out1[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18692), 
          .COUT(n18693), .S0(n1166[5]), .S1(n1166[6]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_7.INIT0 = 16'h5aaa;
    defparam add_183_7.INIT1 = 16'h5aaa;
    defparam add_183_7.INJECT1_0 = "NO";
    defparam add_183_7.INJECT1_1 = "NO";
    CCU2D sub_17_rep_2_add_2_9 (.A0(n2245[7]), .B0(subIn2[7]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[8]), .B1(subIn2[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18757), .COUT(n18758), .S0(n4197), .S1(n4196));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_9.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_9.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_9.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_17_rep_2_add_2_7 (.A0(n2245[5]), .B0(subIn2[5]), .C0(GND_net), 
          .D0(GND_net), .A1(n2245[6]), .B1(subIn2[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18756), .COUT(n18757), .S0(n4199), .S1(n4198));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(228[13:19])
    defparam sub_17_rep_2_add_2_7.INIT0 = 16'h5999;
    defparam sub_17_rep_2_add_2_7.INIT1 = 16'h5999;
    defparam sub_17_rep_2_add_2_7.INJECT1_0 = "NO";
    defparam sub_17_rep_2_add_2_7.INJECT1_1 = "NO";
    CCU2D add_183_5 (.A0(Out1[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18691), 
          .COUT(n18692), .S0(n1166[3]), .S1(n1166[4]));   // c:/users/gebruiker/workspace/lattice/final code software/pid.vhd(315[17:21])
    defparam add_183_5.INIT0 = 16'h5aaa;
    defparam add_183_5.INIT1 = 16'h5aaa;
    defparam add_183_5.INJECT1_0 = "NO";
    defparam add_183_5.INJECT1_1 = "NO";
    
endmodule
