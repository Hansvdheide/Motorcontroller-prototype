// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.9.0.99.2
// Netlist written on Fri Apr 14 12:08:24 2017
//
// Verilog Description of module SPI_loopback_Top
//

module SPI_loopback_Top (CS, SCK, MOSI, MISO, HALL_A_OUT, HALL_B_OUT, 
            HALL_C_OUT, LED1, LED2, LED3, LED4, clkout, H_A_m1, 
            H_B_m1, H_C_m1, MA_m1, MB_m1, MC_m1, H_A_m2, H_B_m2, 
            H_C_m2, MA_m2, MB_m2, MC_m2, H_A_m3, H_B_m3, H_C_m3, 
            MA_m3, MB_m3, MC_m3, H_A_m4, H_B_m4, H_C_m4, MA_m4, 
            MB_m4, MC_m4);   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(24[8:24])
    input CS;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(27[2:4])
    input SCK;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(28[2:5])
    input MOSI;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(29[2:6])
    output MISO;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(30[2:6])
    output HALL_A_OUT;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(33[2:12])
    output HALL_B_OUT;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(34[2:12])
    output HALL_C_OUT;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(35[2:12])
    output LED1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(38[2:6])
    output LED2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(39[2:6])
    output LED3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(40[2:6])
    output LED4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(41[2:6])
    output clkout;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    input H_A_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(47[2:8])
    input H_B_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(48[2:8])
    input H_C_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(49[2:8])
    output [1:0]MA_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(50[2:7])
    output [1:0]MB_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(51[2:7])
    output [1:0]MC_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(52[2:7])
    input H_A_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(55[2:8])
    input H_B_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(56[2:8])
    input H_C_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(57[2:8])
    output [1:0]MA_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(58[2:7])
    output [1:0]MB_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(59[2:7])
    output [1:0]MC_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(60[2:7])
    input H_A_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(63[2:8])
    input H_B_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(64[2:8])
    input H_C_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(65[2:8])
    output [1:0]MA_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(66[2:7])
    output [1:0]MB_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(67[2:7])
    output [1:0]MC_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(68[2:7])
    input H_A_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(71[2:8])
    input H_B_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(72[2:8])
    input H_C_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(73[2:8])
    output [1:0]MA_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(74[2:7])
    output [1:0]MB_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(75[2:7])
    output [1:0]MC_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(76[2:7])
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(88[9:16])
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(30[4:14])
    
    wire GND_net, VCC_net, CS_c, SCK_c, MOSI_c, HALL_A_OUT_c_c, 
        HALL_B_OUT_c_c, HALL_C_OUT_c_c, LED1_c, LED2_c, LED3_c, LED4_c, 
        H_A_m1_c, H_B_m1_c, H_C_m1_c, MA_m1_c_1, MA_m1_c_0, MB_m1_c_1, 
        MB_m1_c_0, MC_m1_c_1, MC_m1_c_0, H_A_m2_c, H_B_m2_c, H_C_m2_c, 
        MA_m2_c_1, MA_m2_c_0, MB_m2_c_1, MB_m2_c_0, MC_m2_c_1, MC_m2_c_0, 
        H_A_m3_c, H_B_m3_c, H_C_m3_c, MA_m3_c_1, MA_m3_c_0, MB_m3_c_1, 
        MB_m3_c_0, MC_m3_c_1, MC_m3_c_0, MA_m4_c_1, MA_m4_c_0, MB_m4_c_1, 
        MB_m4_c_0, MC_m4_c_1, MC_m4_c_0, rst, enable_m1, enable_m2, 
        enable_m3, enable_m4;
    wire [20:0]speed_set_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(99[9:21])
    wire [20:0]speed_set_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(100[9:21])
    wire [20:0]speed_set_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(101[9:21])
    wire [20:0]speed_set_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(102[9:21])
    wire [20:0]speed_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(104[9:17])
    wire [20:0]speed_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(105[9:17])
    wire [20:0]speed_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(106[9:17])
    wire [20:0]speed_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(107[9:17])
    wire [2:0]hallsense_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(110[9:21])
    wire [2:0]hallsense_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(111[9:21])
    wire [2:0]hallsense_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(112[9:21])
    wire [2:0]hallsense_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(113[9:21])
    
    wire PWM_m1, PWM_m2, PWM_m3, PWM_m4;
    wire [9:0]PWMdut_m1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(120[9:18])
    wire [9:0]PWMdut_m2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(121[9:18])
    wire [9:0]PWMdut_m3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(122[9:18])
    wire [9:0]PWMdut_m4;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(123[9:18])
    
    wire dir_m1, dir_m2, dir_m3, dir_m4;
    wire [13:0]start_cnt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(135[9:18])
    
    wire free_m1, free_m2, free_m3, free_m4;
    wire [95:0]send_buffer;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(67[10:21])
    
    wire n3081, n3139, n3057, n3045, n3009, n2951, n19654, n2927, 
        n2915, n2963, n2879, n2821, n2797, n2785, n20183;
    wire [95:0]send_buffer_95__N_346;
    
    wire clkout_c_enable_164, MISO_N_624, n3175, n19650, clkout_c_enable_176, 
        n21544, n18583, n18582, n18581, n18580, n18579, n18578, 
        n18577, n18797, n4132, n18796, n18733, n2833, n3093, n3187, 
        n3211, n3269, n3223, n4883, n62, n63, n64, n65, n66, 
        n67, n68, n69, n70, n71, n72, n73, n74, n75, n10081, 
        n3, clkout_c_enable_257, n7, n5, n19662, n21507, n6, n21598, 
        n21596, n21595, n21593, n21592, n21591, n21590, n21589, 
        n21587, n21585, n22198, n21575, n21574, n21573, n21570, 
        n19656, n22203, n21556, n21555;
    
    VHI i2 (.Z(VCC_net));
    OSCH OSCInst0 (.STDBY(GND_net), .OSC(clkout_c)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCInst0.NOM_FREQ = "38.00";
    OB MA_m2_pad_0 (.I(MA_m2_c_0), .O(MA_m2[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(58[2:7])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    OB HALL_B_OUT_pad (.I(HALL_B_OUT_c_c), .O(HALL_B_OUT));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(34[2:12])
    OB HALL_A_OUT_pad (.I(HALL_A_OUT_c_c), .O(HALL_A_OUT));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(33[2:12])
    OB MA_m2_pad_1 (.I(MA_m2_c_1), .O(MA_m2[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(58[2:7])
    IB H_B_m1_pad (.I(H_B_m1), .O(H_B_m1_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(48[2:8])
    OBZ n4882_pad (.I(MISO_N_624), .T(n4883), .O(MISO));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(64[1] 216[13])
    IB H_A_m1_pad (.I(H_A_m1), .O(H_A_m1_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(47[2:8])
    IB MOSI_pad (.I(MOSI), .O(MOSI_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(29[2:6])
    IB SCK_pad (.I(SCK), .O(SCK_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(28[2:5])
    IB CS_pad (.I(CS), .O(CS_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(27[2:4])
    OB MC_m4_pad_0 (.I(MC_m4_c_0), .O(MC_m4[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(76[2:7])
    OB MC_m4_pad_1 (.I(MC_m4_c_1), .O(MC_m4[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(76[2:7])
    OB MB_m4_pad_0 (.I(MB_m4_c_0), .O(MB_m4[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(75[2:7])
    OB MB_m4_pad_1 (.I(MB_m4_c_1), .O(MB_m4[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(75[2:7])
    OB MC_m1_pad_0 (.I(MC_m1_c_0), .O(MC_m1[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(52[2:7])
    OB MC_m1_pad_1 (.I(MC_m1_c_1), .O(MC_m1[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(52[2:7])
    OB MA_m4_pad_0 (.I(MA_m4_c_0), .O(MA_m4[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_0 (.I(MB_m1_c_0), .O(MB_m1[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(51[2:7])
    OB MA_m4_pad_1 (.I(MA_m4_c_1), .O(MA_m4[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_1 (.I(MB_m1_c_1), .O(MB_m1[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(51[2:7])
    OB MC_m3_pad_0 (.I(MC_m3_c_0), .O(MC_m3[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(68[2:7])
    IB HALL_C_OUT_c_pad (.I(H_C_m4), .O(HALL_C_OUT_c_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(73[2:8])
    OB MA_m1_pad_0 (.I(MA_m1_c_0), .O(MA_m1[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(50[2:7])
    OB MC_m3_pad_1 (.I(MC_m3_c_1), .O(MC_m3[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(68[2:7])
    IB HALL_B_OUT_c_pad (.I(H_B_m4), .O(HALL_B_OUT_c_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(72[2:8])
    OB MA_m1_pad_1 (.I(MA_m1_c_1), .O(MA_m1[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(50[2:7])
    OB MB_m3_pad_0 (.I(MB_m3_c_0), .O(MB_m3[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(67[2:7])
    IB HALL_A_OUT_c_pad (.I(H_A_m4), .O(HALL_A_OUT_c_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(71[2:8])
    OB clkout_pad (.I(clkout_c), .O(clkout));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    OB MB_m3_pad_1 (.I(MB_m3_c_1), .O(MB_m3[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(67[2:7])
    IB H_C_m3_pad (.I(H_C_m3), .O(H_C_m3_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(65[2:8])
    OB LED4_pad (.I(LED4_c), .O(LED4));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(41[2:6])
    OB MA_m3_pad_0 (.I(MA_m3_c_0), .O(MA_m3[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(66[2:7])
    IB H_B_m3_pad (.I(H_B_m3), .O(H_B_m3_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(64[2:8])
    OB LED3_pad (.I(LED3_c), .O(LED3));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(40[2:6])
    OB MA_m3_pad_1 (.I(MA_m3_c_1), .O(MA_m3[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(66[2:7])
    IB H_A_m3_pad (.I(H_A_m3), .O(H_A_m3_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(63[2:8])
    OB LED2_pad (.I(LED2_c), .O(LED2));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(39[2:6])
    OB MC_m2_pad_0 (.I(MC_m2_c_0), .O(MC_m2[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(60[2:7])
    IB H_C_m2_pad (.I(H_C_m2), .O(H_C_m2_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(57[2:8])
    OB LED1_pad (.I(LED1_c), .O(LED1));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(38[2:6])
    OB MC_m2_pad_1 (.I(MC_m2_c_1), .O(MC_m2[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(60[2:7])
    IB H_B_m2_pad (.I(H_B_m2), .O(H_B_m2_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(56[2:8])
    OB HALL_C_OUT_pad (.I(HALL_C_OUT_c_c), .O(HALL_C_OUT));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(35[2:12])
    OB MB_m2_pad_0 (.I(MB_m2_c_0), .O(MB_m2[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(59[2:7])
    IB H_A_m2_pad (.I(H_A_m2), .O(H_A_m2_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(55[2:8])
    OB MB_m2_pad_1 (.I(MB_m2_c_1), .O(MB_m2[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(59[2:7])
    IB H_C_m1_pad (.I(H_C_m1), .O(H_C_m1_c));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(49[2:8])
    FD1P3AX start_cnt_2058__i0 (.D(n75), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i0.GSR = "DISABLED";
    FD1S3AX rst_12 (.D(n21507), .CK(clkout_c), .Q(rst));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_12.GSR = "DISABLED";
    GSR GSR_INST (.GSR(n22203));
    LUT4 i2268_4_lut_rep_298 (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18733), .Z(n21507)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2268_4_lut_rep_298.init = 16'hccc8;
    LUT4 i8944_1_lut_4_lut (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18733), .Z(clkout_c_enable_257)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i8944_1_lut_4_lut.init = 16'h3337;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2D start_cnt_2058_add_4_5 (.A0(start_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18578), .COUT(n18579), .S0(n72), .S1(n71));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_5.INIT0 = 16'hfaaa;
    defparam start_cnt_2058_add_4_5.INIT1 = 16'hfaaa;
    defparam start_cnt_2058_add_4_5.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_5.INJECT1_1 = "NO";
    CCU2D start_cnt_2058_add_4_3 (.A0(start_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18577), .COUT(n18578), .S0(n74), .S1(n73));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_3.INIT0 = 16'hfaaa;
    defparam start_cnt_2058_add_4_3.INIT1 = 16'hfaaa;
    defparam start_cnt_2058_add_4_3.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_3.INJECT1_1 = "NO";
    LUT4 i1745_3_lut_rep_376 (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .Z(n21585)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(128[9:15])
    defparam i1745_3_lut_rep_376.init = 16'h4242;
    LUT4 i17984_2_lut_4_lut (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .D(free_m4), .Z(n3269)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(128[9:15])
    defparam i17984_2_lut_4_lut.init = 16'hffbd;
    CCU2D start_cnt_2058_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18577), .S1(n75));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_1.INIT0 = 16'hF000;
    defparam start_cnt_2058_add_4_1.INIT1 = 16'h0555;
    defparam start_cnt_2058_add_4_1.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(send_buffer[94]), .B(speed_m1[19]), .C(n21555), 
         .D(n21556), .Z(send_buffer_95__N_346[94])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(73[10:15])
    defparam i1_2_lut_4_lut.init = 16'h00ca;
    LUT4 i13580_4_lut (.A(n4132), .B(speed_m3[19]), .C(n21544), .D(speed_m4[19]), 
         .Z(n3)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i13580_4_lut.init = 16'hcac0;
    LUT4 i1653_3_lut_rep_381 (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .Z(n21590)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(127[9:15])
    defparam i1653_3_lut_rep_381.init = 16'h4242;
    LUT4 i17957_2_lut_4_lut (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .D(free_m3), .Z(n3139)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(127[9:15])
    defparam i17957_2_lut_4_lut.init = 16'hffbd;
    LUT4 m1_lut (.Z(n22198)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    LUT4 i7783_2_lut (.A(n21507), .B(n62), .Z(n10081)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam i7783_2_lut.init = 16'heeee;
    LUT4 i1561_3_lut_rep_386 (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .Z(n21595)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(126[9:15])
    defparam i1561_3_lut_rep_386.init = 16'h4242;
    LUT4 i17986_2_lut_4_lut (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .D(free_m2), .Z(n3009)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(126[9:15])
    defparam i17986_2_lut_4_lut.init = 16'hffbd;
    FD1S3AX rst_12_rep_408 (.D(n21507), .CK(clkout_c), .Q(clkout_c_enable_176));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_12_rep_408.GSR = "DISABLED";
    FD1S3AX rst_12_rep_407 (.D(n21507), .CK(clkout_c), .Q(clkout_c_enable_164));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_12_rep_407.GSR = "DISABLED";
    FD1S3AX rst_12_rep_406 (.D(n21507), .CK(clkout_c), .Q(n22203));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(354[3] 361[10])
    defparam rst_12_rep_406.GSR = "DISABLED";
    PFUMX i13584 (.BLUT(n3), .ALUT(n5), .C0(n20183), .Z(n7));
    CCU2D start_cnt_2058_add_4_15 (.A0(start_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18583), .S0(n62));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_15.INIT0 = 16'hfaaa;
    defparam start_cnt_2058_add_4_15.INIT1 = 16'h0000;
    defparam start_cnt_2058_add_4_15.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_15.INJECT1_1 = "NO";
    CCU2D start_cnt_2058_add_4_13 (.A0(start_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18582), .COUT(n18583), .S0(n64), .S1(n63));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_13.INIT0 = 16'hfaaa;
    defparam start_cnt_2058_add_4_13.INIT1 = 16'hfaaa;
    defparam start_cnt_2058_add_4_13.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_13.INJECT1_1 = "NO";
    COMMUTATION_U6 COM_I_M3 (.MB_m3_c_0(MB_m3_c_0), .clkout_c(clkout_c), 
            .MC_m3_c_0(MC_m3_c_0), .MA_m3_c_0(MA_m3_c_0), .LED3_c(LED3_c), 
            .enable_m3(enable_m3), .n3045(n3045), .n21593(n21593), .PWM_m3(PWM_m3), 
            .n3081(n3081), .n21591(n21591), .n19650(n19650), .n21590(n21590), 
            .free_m3(free_m3), .MA_m3_c_1(MA_m3_c_1), .n3139(n3139), .MC_m3_c_1(MC_m3_c_1), 
            .n3093(n3093), .MB_m3_c_1(MB_m3_c_1), .n3057(n3057));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(325[13:24])
    COMMUTATION_U7 COM_I_M2 (.MB_m2_c_0(MB_m2_c_0), .clkout_c(clkout_c), 
            .MC_m2_c_0(MC_m2_c_0), .MA_m2_c_0(MA_m2_c_0), .LED2_c(LED2_c), 
            .enable_m2(enable_m2), .n2915(n2915), .n21598(n21598), .PWM_m2(PWM_m2), 
            .n2951(n2951), .n21596(n21596), .n19656(n19656), .n21595(n21595), 
            .free_m2(free_m2), .MA_m2_c_1(MA_m2_c_1), .n3009(n3009), .MC_m2_c_1(MC_m2_c_1), 
            .n2963(n2963), .MB_m2_c_1(MB_m2_c_1), .n2927(n2927));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(315[13:24])
    COMMUTATION_U8 COM_I_M1 (.MB_m1_c_0(MB_m1_c_0), .clkout_c(clkout_c), 
            .MC_m1_c_0(MC_m1_c_0), .MA_m1_c_0(MA_m1_c_0), .LED1_c(LED1_c), 
            .MA_m1_c_1(MA_m1_c_1), .n19654(n19654), .n2879(n2879), .MC_m1_c_1(MC_m1_c_1), 
            .n2833(n2833), .n2821(n2821), .MB_m1_c_1(MB_m1_c_1), .n2797(n2797), 
            .n2785(n2785), .enable_m1(enable_m1), .n21575(n21575), .PWM_m1(PWM_m1), 
            .n21573(n21573), .n21570(n21570), .free_m1(free_m1));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(305[13:24])
    CCU2D start_cnt_2058_add_4_11 (.A0(start_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18581), .COUT(n18582), .S0(n66), .S1(n65));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_11.INIT0 = 16'hfaaa;
    defparam start_cnt_2058_add_4_11.INIT1 = 16'hfaaa;
    defparam start_cnt_2058_add_4_11.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_11.INJECT1_1 = "NO";
    LUT4 i1469_3_lut_rep_361 (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .Z(n21570)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(125[9:15])
    defparam i1469_3_lut_rep_361.init = 16'h4242;
    LUT4 i17988_2_lut_4_lut (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .D(free_m1), .Z(n2879)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(125[9:15])
    defparam i17988_2_lut_4_lut.init = 16'hffbd;
    SPI SPI_I (.MISO_N_624(MISO_N_624), .clkout_c(clkout_c), .enable_m4(enable_m4), 
        .clkout_c_enable_164(clkout_c_enable_164), .speed_set_m4({speed_set_m4}), 
        .\speed_m4[10] (speed_m4[10]), .CS_c(CS_c), .SCK_c(SCK_c), .enable_m1(enable_m1), 
        .enable_m2(enable_m2), .enable_m3(enable_m3), .\speed_m4[17] (speed_m4[17]), 
        .\speed_m4[18] (speed_m4[18]), .\speed_m4[19] (speed_m4[19]), .\speed_m3[0] (speed_m3[0]), 
        .\speed_m3[1] (speed_m3[1]), .\speed_m3[2] (speed_m3[2]), .\speed_m3[3] (speed_m3[3]), 
        .\speed_m3[4] (speed_m3[4]), .MOSI_c(MOSI_c), .\speed_m3[5] (speed_m3[5]), 
        .\speed_m3[6] (speed_m3[6]), .\speed_m3[7] (speed_m3[7]), .\speed_m3[8] (speed_m3[8]), 
        .\speed_m3[9] (speed_m3[9]), .n21555(n21555), .\speed_m3[10] (speed_m3[10]), 
        .\speed_m3[11] (speed_m3[11]), .\speed_m3[12] (speed_m3[12]), .\speed_m3[13] (speed_m3[13]), 
        .\speed_m3[14] (speed_m3[14]), .\speed_m3[15] (speed_m3[15]), .\speed_m3[16] (speed_m3[16]), 
        .\speed_m3[17] (speed_m3[17]), .\speed_m3[18] (speed_m3[18]), .\speed_m3[19] (speed_m3[19]), 
        .\speed_m2[0] (speed_m2[0]), .\speed_m2[1] (speed_m2[1]), .\speed_m2[2] (speed_m2[2]), 
        .\speed_m2[3] (speed_m2[3]), .\speed_m2[4] (speed_m2[4]), .\speed_m2[5] (speed_m2[5]), 
        .\speed_m4[5] (speed_m4[5]), .\speed_m4[4] (speed_m4[4]), .\speed_m2[6] (speed_m2[6]), 
        .\speed_m2[7] (speed_m2[7]), .\speed_m2[8] (speed_m2[8]), .\speed_m2[9] (speed_m2[9]), 
        .\speed_m2[10] (speed_m2[10]), .\speed_m2[11] (speed_m2[11]), .\speed_m2[12] (speed_m2[12]), 
        .\speed_m2[13] (speed_m2[13]), .\speed_m2[14] (speed_m2[14]), .\speed_m2[15] (speed_m2[15]), 
        .\speed_m2[16] (speed_m2[16]), .\speed_m2[17] (speed_m2[17]), .\speed_m2[18] (speed_m2[18]), 
        .\speed_m2[19] (speed_m2[19]), .\speed_m1[0] (speed_m1[0]), .\speed_m1[1] (speed_m1[1]), 
        .\speed_m1[2] (speed_m1[2]), .\speed_m1[3] (speed_m1[3]), .\speed_m1[4] (speed_m1[4]), 
        .\speed_m4[7] (speed_m4[7]), .\speed_m4[6] (speed_m4[6]), .\speed_m1[5] (speed_m1[5]), 
        .\speed_m1[6] (speed_m1[6]), .\speed_m1[7] (speed_m1[7]), .\speed_m1[8] (speed_m1[8]), 
        .\speed_m1[9] (speed_m1[9]), .\speed_m1[10] (speed_m1[10]), .\speed_m1[11] (speed_m1[11]), 
        .\speed_m1[12] (speed_m1[12]), .\speed_m1[13] (speed_m1[13]), .\speed_m1[14] (speed_m1[14]), 
        .\speed_m1[15] (speed_m1[15]), .\speed_m1[16] (speed_m1[16]), .\speed_m1[17] (speed_m1[17]), 
        .\speed_m1[18] (speed_m1[18]), .\speed_m4[8] (speed_m4[8]), .\send_buffer[94] (send_buffer[94]), 
        .\speed_m1[19] (speed_m1[19]), .\speed_m4[0] (speed_m4[0]), .\speed_m4[1] (speed_m4[1]), 
        .\speed_m4[2] (speed_m4[2]), .\speed_m4[3] (speed_m4[3]), .speed_set_m3({speed_set_m3}), 
        .speed_set_m2({speed_set_m2}), .speed_set_m1({speed_set_m1}), .free_m4(free_m4), 
        .hallsense_m4({hallsense_m4}), .n19662(n19662), .n22203(n22203), 
        .\speed_m4[12] (speed_m4[12]), .GND_net(GND_net), .clkout_c_enable_176(clkout_c_enable_176), 
        .rst(rst), .\send_buffer_95__N_346[94] (send_buffer_95__N_346[94]), 
        .free_m2(free_m2), .hallsense_m2({hallsense_m2}), .n19656(n19656), 
        .n4883(n4883), .n21556(n21556), .\speed_m4[16] (speed_m4[16]), 
        .dir_m2(dir_m2), .n2915(n2915), .n2951(n2951), .hallsense_m3({hallsense_m3}), 
        .n21592(n21592), .dir_m3(dir_m3), .n3045(n3045), .n3081(n3081), 
        .dir_m4(dir_m4), .n3175(n3175), .n3211(n3211), .hallsense_m1({hallsense_m1}), 
        .n21574(n21574), .dir_m1(dir_m1), .n2785(n2785), .n2821(n2821), 
        .\speed_m4[11] (speed_m4[11]), .\speed_m4[13] (speed_m4[13]), .\speed_m4[14] (speed_m4[14]), 
        .\speed_m4[9] (speed_m4[9]), .\speed_m4[15] (speed_m4[15]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(293[10:13])
    LUT4 i3_4_lut (.A(n18797), .B(start_cnt[10]), .C(start_cnt[9]), .D(start_cnt[8]), 
         .Z(n18733)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    CCU2D start_cnt_2058_add_4_9 (.A0(start_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18580), .COUT(n18581), .S0(n68), .S1(n67));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_9.INIT0 = 16'hfaaa;
    defparam start_cnt_2058_add_4_9.INIT1 = 16'hfaaa;
    defparam start_cnt_2058_add_4_9.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_9.INJECT1_1 = "NO";
    CCU2D start_cnt_2058_add_4_7 (.A0(start_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18579), .COUT(n18580), .S0(n70), .S1(n69));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058_add_4_7.INIT0 = 16'hfaaa;
    defparam start_cnt_2058_add_4_7.INIT1 = 16'hfaaa;
    defparam start_cnt_2058_add_4_7.INJECT1_0 = "NO";
    defparam start_cnt_2058_add_4_7.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_166 (.A(n18796), .B(n6), .C(start_cnt[6]), .D(start_cnt[4]), 
         .Z(n18797)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_166.init = 16'hfefc;
    LUT4 i3_4_lut_adj_167 (.A(start_cnt[0]), .B(start_cnt[3]), .C(start_cnt[2]), 
         .D(start_cnt[1]), .Z(n18796)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_167.init = 16'hfffe;
    LUT4 i2_2_lut (.A(start_cnt[7]), .B(start_cnt[5]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    HALL_U4 HALL_I_M2 (.clk_1mhz(clk_1mhz), .\speed_m2[0] (speed_m2[0]), 
            .hallsense_m2({hallsense_m2}), .clkout_c_enable_176(clkout_c_enable_176), 
            .clkout_c_enable_164(clkout_c_enable_164), .H_C_m2_c(H_C_m2_c), 
            .H_B_m2_c(H_B_m2_c), .H_A_m2_c(H_A_m2_c), .\speed_m2[1] (speed_m2[1]), 
            .\speed_m2[2] (speed_m2[2]), .\speed_m2[3] (speed_m2[3]), .\speed_m2[4] (speed_m2[4]), 
            .\speed_m2[5] (speed_m2[5]), .\speed_m2[6] (speed_m2[6]), .\speed_m2[7] (speed_m2[7]), 
            .\speed_m2[8] (speed_m2[8]), .\speed_m2[9] (speed_m2[9]), .\speed_m2[10] (speed_m2[10]), 
            .\speed_m2[11] (speed_m2[11]), .\speed_m2[12] (speed_m2[12]), 
            .\speed_m2[13] (speed_m2[13]), .\speed_m2[14] (speed_m2[14]), 
            .\speed_m2[15] (speed_m2[15]), .\speed_m2[16] (speed_m2[16]), 
            .\speed_m2[17] (speed_m2[17]), .\speed_m2[18] (speed_m2[18]), 
            .\speed_m2[19] (speed_m2[19]), .GND_net(GND_net), .n22198(n22198));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(312[14:18])
    HALL_U3 HALL_I_M3 (.clk_1mhz(clk_1mhz), .\speed_m3[0] (speed_m3[0]), 
            .hallsense_m3({hallsense_m3}), .clkout_c_enable_176(clkout_c_enable_176), 
            .H_A_m3_c(H_A_m3_c), .H_B_m3_c(H_B_m3_c), .H_C_m3_c(H_C_m3_c), 
            .clkout_c_enable_164(clkout_c_enable_164), .\speed_m3[1] (speed_m3[1]), 
            .\speed_m3[2] (speed_m3[2]), .\speed_m3[3] (speed_m3[3]), .\speed_m3[4] (speed_m3[4]), 
            .\speed_m3[5] (speed_m3[5]), .\speed_m3[6] (speed_m3[6]), .\speed_m3[7] (speed_m3[7]), 
            .\speed_m3[8] (speed_m3[8]), .\speed_m3[9] (speed_m3[9]), .\speed_m3[10] (speed_m3[10]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_m3[12] (speed_m3[12]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_m3[14] (speed_m3[14]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_m3[16] (speed_m3[16]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_m3[18] (speed_m3[18]), 
            .\speed_m3[19] (speed_m3[19]), .GND_net(GND_net), .n22198(n22198));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(322[14:18])
    HALL_U5 HALL_I_M1 (.clk_1mhz(clk_1mhz), .\speed_m1[0] (speed_m1[0]), 
            .hallsense_m1({hallsense_m1}), .clkout_c_enable_164(clkout_c_enable_164), 
            .clkout_c_enable_176(clkout_c_enable_176), .H_A_m1_c(H_A_m1_c), 
            .H_B_m1_c(H_B_m1_c), .H_C_m1_c(H_C_m1_c), .\speed_m1[1] (speed_m1[1]), 
            .\speed_m1[2] (speed_m1[2]), .\speed_m1[3] (speed_m1[3]), .\speed_m1[4] (speed_m1[4]), 
            .\speed_m1[5] (speed_m1[5]), .\speed_m1[6] (speed_m1[6]), .\speed_m1[7] (speed_m1[7]), 
            .\speed_m1[8] (speed_m1[8]), .\speed_m1[9] (speed_m1[9]), .\speed_m1[10] (speed_m1[10]), 
            .\speed_m1[11] (speed_m1[11]), .\speed_m1[12] (speed_m1[12]), 
            .\speed_m1[13] (speed_m1[13]), .\speed_m1[14] (speed_m1[14]), 
            .\speed_m1[15] (speed_m1[15]), .\speed_m1[16] (speed_m1[16]), 
            .\speed_m1[17] (speed_m1[17]), .\speed_m1[18] (speed_m1[18]), 
            .\speed_m1[19] (speed_m1[19]), .GND_net(GND_net), .n22198(n22198));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(302[14:18])
    COMMUTATION COM_I_M4 (.MB_m4_c_0(MB_m4_c_0), .clkout_c(clkout_c), .MC_m4_c_0(MC_m4_c_0), 
            .MA_m4_c_0(MA_m4_c_0), .LED4_c(LED4_c), .enable_m4(enable_m4), 
            .n3175(n3175), .n21589(n21589), .PWM_m4(PWM_m4), .n3211(n3211), 
            .n21587(n21587), .n19662(n19662), .n21585(n21585), .free_m4(free_m4), 
            .MA_m4_c_1(MA_m4_c_1), .n3269(n3269), .MC_m4_c_1(MC_m4_c_1), 
            .n3223(n3223), .MB_m4_c_1(MB_m4_c_1), .n3187(n3187));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(335[13:24])
    CLKDIV CLKDIV_I (.clk_N_683(clk_N_683), .clkout_c(clkout_c), .clk_1mhz(clk_1mhz), 
           .pwm_clk(pwm_clk), .GND_net(GND_net));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(288[14:20])
    PWMGENERATOR_U0 PWM_I_M3 (.PWM_m3(PWM_m3), .pwm_clk(pwm_clk), .free_m3(free_m3), 
            .clkout_c_enable_176(clkout_c_enable_176), .hallsense_m3({hallsense_m3}), 
            .n21591(n21591), .enable_m3(enable_m3), .n3093(n3093), .PWMdut_m3({PWMdut_m3}), 
            .GND_net(GND_net), .n21592(n21592), .n19650(n19650), .n21593(n21593), 
            .n3057(n3057));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(328[13:25])
    PWMGENERATOR_U1 PWM_I_M2 (.PWM_m2(PWM_m2), .pwm_clk(pwm_clk), .free_m2(free_m2), 
            .clkout_c_enable_176(clkout_c_enable_176), .PWMdut_m2({PWMdut_m2}), 
            .GND_net(GND_net), .hallsense_m2({hallsense_m2}), .n21596(n21596), 
            .enable_m2(enable_m2), .n2963(n2963), .n21598(n21598), .n2927(n2927));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(318[13:25])
    PWMGENERATOR_U2 PWM_I_M1 (.GND_net(GND_net), .PWMdut_m1({PWMdut_m1}), 
            .PWM_m1(PWM_m1), .pwm_clk(pwm_clk), .free_m1(free_m1), .clkout_c_enable_164(clkout_c_enable_164), 
            .hallsense_m1({hallsense_m1}), .n21573(n21573), .enable_m1(enable_m1), 
            .n2833(n2833), .n21574(n21574), .n19654(n19654), .n21575(n21575), 
            .n2797(n2797));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(308[13:25])
    \PID(16000000,160000000,10000000)  PID_I (.clk_N_683(clk_N_683), .GND_net(GND_net), 
            .PWMdut_m3({PWMdut_m3}), .dir_m2(dir_m2), .dir_m3(dir_m3), 
            .dir_m1(dir_m1), .dir_m4(dir_m4), .speed_set_m2({speed_set_m2}), 
            .speed_set_m1({speed_set_m1}), .VCC_net(VCC_net), .speed_set_m4({speed_set_m4}), 
            .\speed_m4[0] (speed_m4[0]), .\speed_m3[0] (speed_m3[0]), .n21544(n21544), 
            .n4132(n4132), .\speed_m3[3] (speed_m3[3]), .\speed_m2[3] (speed_m2[3]), 
            .\speed_m4[12] (speed_m4[12]), .\speed_m3[7] (speed_m3[7]), 
            .\speed_m2[7] (speed_m2[7]), .\speed_m3[8] (speed_m3[8]), .\speed_m2[8] (speed_m2[8]), 
            .\speed_m3[9] (speed_m3[9]), .\speed_m2[9] (speed_m2[9]), .\speed_m3[12] (speed_m3[12]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_m4[9] (speed_m4[9]), 
            .\speed_m4[8] (speed_m4[8]), .\speed_m4[18] (speed_m4[18]), 
            .\speed_m3[18] (speed_m3[18]), .\speed_m4[7] (speed_m4[7]), 
            .\speed_m4[3] (speed_m4[3]), .\speed_m4[17] (speed_m4[17]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_m4[16] (speed_m4[16]), 
            .\speed_m3[16] (speed_m3[16]), .\speed_m4[15] (speed_m4[15]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_m4[14] (speed_m4[14]), 
            .\speed_m3[14] (speed_m3[14]), .\speed_m4[13] (speed_m4[13]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_m4[11] (speed_m4[11]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_m4[10] (speed_m4[10]), 
            .\speed_m3[10] (speed_m3[10]), .\speed_m4[6] (speed_m4[6]), 
            .\speed_m3[6] (speed_m3[6]), .\speed_m4[5] (speed_m4[5]), .\speed_m3[5] (speed_m3[5]), 
            .\speed_m4[4] (speed_m4[4]), .\speed_m3[4] (speed_m3[4]), .\speed_m4[2] (speed_m4[2]), 
            .\speed_m3[2] (speed_m3[2]), .n22203(n22203), .\speed_m4[1] (speed_m4[1]), 
            .\speed_m3[1] (speed_m3[1]), .\speed_m1[0] (speed_m1[0]), .\speed_m2[0] (speed_m2[0]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_m2[18] (speed_m2[18]), 
            .\speed_m1[17] (speed_m1[17]), .\speed_m2[17] (speed_m2[17]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_m2[16] (speed_m2[16]), 
            .\speed_m1[15] (speed_m1[15]), .\speed_m2[15] (speed_m2[15]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_m2[14] (speed_m2[14]), 
            .\speed_m1[13] (speed_m1[13]), .\speed_m2[13] (speed_m2[13]), 
            .\speed_m1[11] (speed_m1[11]), .\speed_m2[11] (speed_m2[11]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_m2[10] (speed_m2[10]), 
            .\speed_m1[6] (speed_m1[6]), .\speed_m2[6] (speed_m2[6]), .\speed_m1[5] (speed_m1[5]), 
            .\speed_m2[5] (speed_m2[5]), .\speed_m1[4] (speed_m1[4]), .\speed_m2[4] (speed_m2[4]), 
            .\speed_m1[2] (speed_m1[2]), .\speed_m2[2] (speed_m2[2]), .\speed_m1[1] (speed_m1[1]), 
            .\speed_m2[1] (speed_m2[1]), .\speed_m1[19] (speed_m1[19]), 
            .\speed_m2[19] (speed_m2[19]), .n5(n5), .\speed_m1[12] (speed_m1[12]), 
            .\speed_m1[9] (speed_m1[9]), .\speed_m1[8] (speed_m1[8]), .\speed_m1[7] (speed_m1[7]), 
            .\speed_m1[3] (speed_m1[3]), .PWMdut_m2({PWMdut_m2}), .PWMdut_m1({PWMdut_m1}), 
            .speed_set_m3({speed_set_m3}), .n7(n7), .n20183(n20183), .PWMdut_m4({PWMdut_m4}));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(297[10:13])
    PWMGENERATOR PWM_I_M4 (.PWM_m4(PWM_m4), .pwm_clk(pwm_clk), .free_m4(free_m4), 
            .clkout_c_enable_176(clkout_c_enable_176), .hallsense_m4({hallsense_m4}), 
            .n21587(n21587), .enable_m4(enable_m4), .n3223(n3223), .n21589(n21589), 
            .n3187(n3187), .PWMdut_m4({PWMdut_m4}), .GND_net(GND_net));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(338[13:25])
    HALL HALL_I_M4 (.clk_1mhz(clk_1mhz), .\speed_m4[0] (speed_m4[0]), .clkout_c_enable_176(clkout_c_enable_176), 
         .hallsense_m4({hallsense_m4}), .HALL_A_OUT_c_c(HALL_A_OUT_c_c), 
         .HALL_B_OUT_c_c(HALL_B_OUT_c_c), .HALL_C_OUT_c_c(HALL_C_OUT_c_c), 
         .clkout_c_enable_164(clkout_c_enable_164), .\speed_m4[1] (speed_m4[1]), 
         .\speed_m4[2] (speed_m4[2]), .\speed_m4[3] (speed_m4[3]), .\speed_m4[4] (speed_m4[4]), 
         .\speed_m4[5] (speed_m4[5]), .\speed_m4[6] (speed_m4[6]), .\speed_m4[7] (speed_m4[7]), 
         .\speed_m4[8] (speed_m4[8]), .\speed_m4[9] (speed_m4[9]), .\speed_m4[10] (speed_m4[10]), 
         .\speed_m4[11] (speed_m4[11]), .\speed_m4[12] (speed_m4[12]), .\speed_m4[13] (speed_m4[13]), 
         .\speed_m4[14] (speed_m4[14]), .\speed_m4[15] (speed_m4[15]), .\speed_m4[16] (speed_m4[16]), 
         .\speed_m4[17] (speed_m4[17]), .\speed_m4[18] (speed_m4[18]), .\speed_m4[19] (speed_m4[19]), 
         .GND_net(GND_net), .n22198(n22198));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(332[14:18])
    FD1P3AX start_cnt_2058__i1 (.D(n74), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i1.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i2 (.D(n73), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i2.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i3 (.D(n72), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i3.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i4 (.D(n71), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i4.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i5 (.D(n70), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i5.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i6 (.D(n69), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i6.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i7 (.D(n68), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i7.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i8 (.D(n67), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i8.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i9 (.D(n66), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i9.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i10 (.D(n65), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i10.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i11 (.D(n64), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i11.GSR = "DISABLED";
    FD1P3AX start_cnt_2058__i12 (.D(n63), .SP(clkout_c_enable_257), .CK(clkout_c), 
            .Q(start_cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i12.GSR = "DISABLED";
    FD1S3AX start_cnt_2058__i13 (.D(n10081), .CK(clkout_c), .Q(start_cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(359[18:27])
    defparam start_cnt_2058__i13.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module COMMUTATION_U6
//

module COMMUTATION_U6 (MB_m3_c_0, clkout_c, MC_m3_c_0, MA_m3_c_0, LED3_c, 
            enable_m3, n3045, n21593, PWM_m3, n3081, n21591, n19650, 
            n21590, free_m3, MA_m3_c_1, n3139, MC_m3_c_1, n3093, 
            MB_m3_c_1, n3057);
    output MB_m3_c_0;
    input clkout_c;
    output MC_m3_c_0;
    output MA_m3_c_0;
    output LED3_c;
    input enable_m3;
    input n3045;
    input n21593;
    input PWM_m3;
    input n3081;
    input n21591;
    input n19650;
    input n21590;
    input free_m3;
    output MA_m3_c_1;
    input n3139;
    output MC_m3_c_1;
    input n3093;
    output MB_m3_c_1;
    input n3057;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n18806, n18798, n19651, clkout_c_enable_8;
    
    FD1S3IX MospairB_i1 (.D(n18806), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18798), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19651), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_8), .CK(clkout_c), 
            .Q(LED3_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10095_1_lut (.A(enable_m3), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i10095_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3045), .B(n21593), .C(PWM_m3), .Z(n18806)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_165 (.A(n3081), .B(n21591), .C(PWM_m3), .Z(n18798)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_165.init = 16'hbfbf;
    LUT4 i17847_3_lut (.A(n19650), .B(PWM_m3), .C(n21590), .Z(n19651)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17847_3_lut.init = 16'hbfbf;
    LUT4 i17965_2_lut (.A(free_m3), .B(enable_m3), .Z(clkout_c_enable_8)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i17965_2_lut.init = 16'h7777;
    FD1S3IX MospairA_i2 (.D(n3139), .CK(clkout_c), .CD(n19650), .Q(MA_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3081), .CK(clkout_c), .CD(n3093), .Q(MC_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3045), .CK(clkout_c), .CD(n3057), .Q(MB_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION_U7
//

module COMMUTATION_U7 (MB_m2_c_0, clkout_c, MC_m2_c_0, MA_m2_c_0, LED2_c, 
            enable_m2, n2915, n21598, PWM_m2, n2951, n21596, n19656, 
            n21595, free_m2, MA_m2_c_1, n3009, MC_m2_c_1, n2963, 
            MB_m2_c_1, n2927);
    output MB_m2_c_0;
    input clkout_c;
    output MC_m2_c_0;
    output MA_m2_c_0;
    output LED2_c;
    input enable_m2;
    input n2915;
    input n21598;
    input PWM_m2;
    input n2951;
    input n21596;
    input n19656;
    input n21595;
    input free_m2;
    output MA_m2_c_1;
    input n3009;
    output MC_m2_c_1;
    input n2963;
    output MB_m2_c_1;
    input n2927;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n18808, n18807, n19657, clkout_c_enable_5;
    
    FD1S3IX MospairB_i1 (.D(n18808), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18807), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19657), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_5), .CK(clkout_c), 
            .Q(LED2_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10094_1_lut (.A(enable_m2), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i10094_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2915), .B(n21598), .C(PWM_m2), .Z(n18808)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_164 (.A(n2951), .B(n21596), .C(PWM_m2), .Z(n18807)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_164.init = 16'hbfbf;
    LUT4 i17912_3_lut (.A(n19656), .B(PWM_m2), .C(n21595), .Z(n19657)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17912_3_lut.init = 16'hbfbf;
    LUT4 i17968_2_lut (.A(free_m2), .B(enable_m2), .Z(clkout_c_enable_5)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i17968_2_lut.init = 16'h7777;
    FD1S3IX MospairA_i2 (.D(n3009), .CK(clkout_c), .CD(n19656), .Q(MA_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n2951), .CK(clkout_c), .CD(n2963), .Q(MC_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2915), .CK(clkout_c), .CD(n2927), .Q(MB_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=315, LSE_RLINE=315 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION_U8
//

module COMMUTATION_U8 (MB_m1_c_0, clkout_c, MC_m1_c_0, MA_m1_c_0, LED1_c, 
            MA_m1_c_1, n19654, n2879, MC_m1_c_1, n2833, n2821, MB_m1_c_1, 
            n2797, n2785, enable_m1, n21575, PWM_m1, n21573, n21570, 
            free_m1);
    output MB_m1_c_0;
    input clkout_c;
    output MC_m1_c_0;
    output MA_m1_c_0;
    output LED1_c;
    output MA_m1_c_1;
    input n19654;
    input n2879;
    output MC_m1_c_1;
    input n2833;
    input n2821;
    output MB_m1_c_1;
    input n2797;
    input n2785;
    input enable_m1;
    input n21575;
    input PWM_m1;
    input n21573;
    input n21570;
    input free_m1;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n18810, n18809, n19655, clkout_c_enable_4;
    
    FD1S3IX MospairB_i1 (.D(n18810), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18809), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19655), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_4), .CK(clkout_c), 
            .Q(LED1_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    FD1S3IX MospairA_i2 (.D(n2879), .CK(clkout_c), .CD(n19654), .Q(MA_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n2821), .CK(clkout_c), .CD(n2833), .Q(MC_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2785), .CK(clkout_c), .CD(n2797), .Q(MB_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=305, LSE_RLINE=305 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i10093_1_lut (.A(enable_m1), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i10093_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2785), .B(n21575), .C(PWM_m1), .Z(n18810)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_163 (.A(n2821), .B(n21573), .C(PWM_m1), .Z(n18809)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_163.init = 16'hbfbf;
    LUT4 i17915_3_lut (.A(n19654), .B(PWM_m1), .C(n21570), .Z(n19655)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17915_3_lut.init = 16'hbfbf;
    LUT4 i17971_2_lut (.A(free_m1), .B(enable_m1), .Z(clkout_c_enable_4)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i17971_2_lut.init = 16'h7777;
    
endmodule
//
// Verilog Description of module SPI
//

module SPI (MISO_N_624, clkout_c, enable_m4, clkout_c_enable_164, speed_set_m4, 
            \speed_m4[10] , CS_c, SCK_c, enable_m1, enable_m2, enable_m3, 
            \speed_m4[17] , \speed_m4[18] , \speed_m4[19] , \speed_m3[0] , 
            \speed_m3[1] , \speed_m3[2] , \speed_m3[3] , \speed_m3[4] , 
            MOSI_c, \speed_m3[5] , \speed_m3[6] , \speed_m3[7] , \speed_m3[8] , 
            \speed_m3[9] , n21555, \speed_m3[10] , \speed_m3[11] , \speed_m3[12] , 
            \speed_m3[13] , \speed_m3[14] , \speed_m3[15] , \speed_m3[16] , 
            \speed_m3[17] , \speed_m3[18] , \speed_m3[19] , \speed_m2[0] , 
            \speed_m2[1] , \speed_m2[2] , \speed_m2[3] , \speed_m2[4] , 
            \speed_m2[5] , \speed_m4[5] , \speed_m4[4] , \speed_m2[6] , 
            \speed_m2[7] , \speed_m2[8] , \speed_m2[9] , \speed_m2[10] , 
            \speed_m2[11] , \speed_m2[12] , \speed_m2[13] , \speed_m2[14] , 
            \speed_m2[15] , \speed_m2[16] , \speed_m2[17] , \speed_m2[18] , 
            \speed_m2[19] , \speed_m1[0] , \speed_m1[1] , \speed_m1[2] , 
            \speed_m1[3] , \speed_m1[4] , \speed_m4[7] , \speed_m4[6] , 
            \speed_m1[5] , \speed_m1[6] , \speed_m1[7] , \speed_m1[8] , 
            \speed_m1[9] , \speed_m1[10] , \speed_m1[11] , \speed_m1[12] , 
            \speed_m1[13] , \speed_m1[14] , \speed_m1[15] , \speed_m1[16] , 
            \speed_m1[17] , \speed_m1[18] , \speed_m4[8] , \send_buffer[94] , 
            \speed_m1[19] , \speed_m4[0] , \speed_m4[1] , \speed_m4[2] , 
            \speed_m4[3] , speed_set_m3, speed_set_m2, speed_set_m1, 
            free_m4, hallsense_m4, n19662, n22203, \speed_m4[12] , 
            GND_net, clkout_c_enable_176, rst, \send_buffer_95__N_346[94] , 
            free_m2, hallsense_m2, n19656, n4883, n21556, \speed_m4[16] , 
            dir_m2, n2915, n2951, hallsense_m3, n21592, dir_m3, 
            n3045, n3081, dir_m4, n3175, n3211, hallsense_m1, n21574, 
            dir_m1, n2785, n2821, \speed_m4[11] , \speed_m4[13] , 
            \speed_m4[14] , \speed_m4[9] , \speed_m4[15] );
    output MISO_N_624;
    input clkout_c;
    output enable_m4;
    input clkout_c_enable_164;
    output [20:0]speed_set_m4;
    input \speed_m4[10] ;
    input CS_c;
    input SCK_c;
    output enable_m1;
    output enable_m2;
    output enable_m3;
    input \speed_m4[17] ;
    input \speed_m4[18] ;
    input \speed_m4[19] ;
    input \speed_m3[0] ;
    input \speed_m3[1] ;
    input \speed_m3[2] ;
    input \speed_m3[3] ;
    input \speed_m3[4] ;
    input MOSI_c;
    input \speed_m3[5] ;
    input \speed_m3[6] ;
    input \speed_m3[7] ;
    input \speed_m3[8] ;
    input \speed_m3[9] ;
    output n21555;
    input \speed_m3[10] ;
    input \speed_m3[11] ;
    input \speed_m3[12] ;
    input \speed_m3[13] ;
    input \speed_m3[14] ;
    input \speed_m3[15] ;
    input \speed_m3[16] ;
    input \speed_m3[17] ;
    input \speed_m3[18] ;
    input \speed_m3[19] ;
    input \speed_m2[0] ;
    input \speed_m2[1] ;
    input \speed_m2[2] ;
    input \speed_m2[3] ;
    input \speed_m2[4] ;
    input \speed_m2[5] ;
    input \speed_m4[5] ;
    input \speed_m4[4] ;
    input \speed_m2[6] ;
    input \speed_m2[7] ;
    input \speed_m2[8] ;
    input \speed_m2[9] ;
    input \speed_m2[10] ;
    input \speed_m2[11] ;
    input \speed_m2[12] ;
    input \speed_m2[13] ;
    input \speed_m2[14] ;
    input \speed_m2[15] ;
    input \speed_m2[16] ;
    input \speed_m2[17] ;
    input \speed_m2[18] ;
    input \speed_m2[19] ;
    input \speed_m1[0] ;
    input \speed_m1[1] ;
    input \speed_m1[2] ;
    input \speed_m1[3] ;
    input \speed_m1[4] ;
    input \speed_m4[7] ;
    input \speed_m4[6] ;
    input \speed_m1[5] ;
    input \speed_m1[6] ;
    input \speed_m1[7] ;
    input \speed_m1[8] ;
    input \speed_m1[9] ;
    input \speed_m1[10] ;
    input \speed_m1[11] ;
    input \speed_m1[12] ;
    input \speed_m1[13] ;
    input \speed_m1[14] ;
    input \speed_m1[15] ;
    input \speed_m1[16] ;
    input \speed_m1[17] ;
    input \speed_m1[18] ;
    input \speed_m4[8] ;
    output \send_buffer[94] ;
    input \speed_m1[19] ;
    input \speed_m4[0] ;
    input \speed_m4[1] ;
    input \speed_m4[2] ;
    input \speed_m4[3] ;
    output [20:0]speed_set_m3;
    output [20:0]speed_set_m2;
    output [20:0]speed_set_m1;
    input free_m4;
    input [2:0]hallsense_m4;
    output n19662;
    input n22203;
    input \speed_m4[12] ;
    input GND_net;
    input clkout_c_enable_176;
    input rst;
    input \send_buffer_95__N_346[94] ;
    input free_m2;
    input [2:0]hallsense_m2;
    output n19656;
    output n4883;
    output n21556;
    input \speed_m4[16] ;
    input dir_m2;
    output n2915;
    output n2951;
    input [2:0]hallsense_m3;
    input n21592;
    input dir_m3;
    output n3045;
    output n3081;
    input dir_m4;
    output n3175;
    output n3211;
    input [2:0]hallsense_m1;
    input n21574;
    input dir_m1;
    output n2785;
    output n2821;
    input \speed_m4[11] ;
    input \speed_m4[13] ;
    input \speed_m4[14] ;
    input \speed_m4[9] ;
    input \speed_m4[15] ;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    
    wire MISO_N_670, enable_m1_N_633, enable_m4_N_649, CSold, n22201, 
        SCKold, SCKlatched, clkout_c_enable_245, n12557;
    wire [83:0]n169;
    wire [95:0]send_buffer;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(67[10:21])
    
    wire n22202;
    wire [95:0]MISOb_N_666;
    
    wire CSlatched, clkout_c_enable_61;
    wire [95:0]recv_buffer;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(68[10:21])
    
    wire enable_m1_N_627, enable_m2_N_635, enable_m3_N_642, MISO_N_625, 
        n21581, MISOb, MISOb_N_660, n21481, n21580, n21480, n21525;
    wire [95:0]send_buffer_95__N_346;
    
    wire clkout_c_enable_96, n12577, n12597, n12617, n3479, n3455, 
        n39_adj_1886, n40_adj_1887, n36_adj_1888, n28_adj_1889, n38_adj_1890, 
        n32_adj_1891, n21588, n34_adj_1892, n24_adj_1893, n18634, 
        n3431, n18633, n18632, n18631, n18630, n18629, n18628, 
        n18627, n3383, n18626, n21597, n18625, n18624, n18623, 
        n18622, n18621, n18620, n3359, n18619, n18618, n18617, 
        n18616, n18615, n18614, n18613, n18612, n18611, n18610, 
        n3335, n18609, n18608, n18607, n18606, n18605, n18604, 
        n18603, n3407, n18602, n18601, n18600, n18599, n18598, 
        n18597, n18596, n18595, n18662, n18594, n18661, n18660, 
        n18659, n18658, n18657, n18656, n18655, n18654, n18653, 
        n3311, n39_adj_1894, n40_adj_1895, n36_adj_1896, n28_adj_1897, 
        n38_adj_1898, n32_adj_1899, n34_adj_1900, n24_adj_1901, n18652, 
        n18651, n18650, n18649, n18648, n18647, n18646, n18727, 
        n18726, n18725, n18724, n18723, n18722, n39_adj_1902, n40_adj_1903, 
        n36_adj_1904, n28_adj_1905, n38_adj_1906, n32_adj_1907, n34_adj_1908, 
        n24_adj_1909, n39_adj_1910, n40_adj_1911, n36_adj_1912, n28_adj_1913, 
        n38_adj_1914, n32_adj_1915, n34_adj_1916, n24_adj_1917, n18721, 
        n18720, n18719, n18718;
    
    FD1S3AX MISO_124 (.D(MISO_N_670), .CK(clkout_c), .Q(MISO_N_624)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISO_124.GSR = "DISABLED";
    FD1P3AX enable_m4_112 (.D(enable_m4_N_649), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m4));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m4_112.GSR = "ENABLED";
    FD1P3AX CSold_113 (.D(n22201), .SP(clkout_c_enable_164), .CK(clkout_c), 
            .Q(CSold));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_113.GSR = "DISABLED";
    FD1P3AX SCKold_114 (.D(SCKlatched), .SP(clkout_c_enable_164), .CK(clkout_c), 
            .Q(SCKold));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKold_114.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i0 (.D(n169[0]), .SP(clkout_c_enable_245), .PD(n12557), 
            .CK(clkout_c), .Q(speed_set_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i0.GSR = "DISABLED";
    LUT4 mux_9_i23_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[22]), .C(\speed_m4[10] ), 
         .D(n22202), .Z(MISOb_N_666[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX CSlatched_115 (.D(CS_c), .SP(clkout_c_enable_164), .CK(clkout_c), 
            .Q(CSlatched));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_115.GSR = "DISABLED";
    FD1P3AX SCKlatched_116 (.D(SCK_c), .SP(clkout_c_enable_164), .CK(clkout_c), 
            .Q(SCKlatched));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKlatched_116.GSR = "DISABLED";
    FD1P3AX \SPI__7_rep_4__i0  (.D(recv_buffer[13]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(n169[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7_rep_4__i0 .GSR = "DISABLED";
    FD1P3AX enable_m1_109 (.D(enable_m1_N_627), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m1));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m1_109.GSR = "ENABLED";
    FD1P3AX enable_m2_110 (.D(enable_m2_N_635), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m2));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m2_110.GSR = "ENABLED";
    FD1P3AX enable_m3_111 (.D(enable_m3_N_642), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m3));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m3_111.GSR = "ENABLED";
    FD1P3AX i101_125 (.D(n21581), .SP(clkout_c_enable_164), .CK(clkout_c), 
            .Q(MISO_N_625));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i101_125.GSR = "DISABLED";
    FD1P3AX MISOb_118 (.D(MISOb_N_660), .SP(clkout_c_enable_164), .CK(clkout_c), 
            .Q(MISOb));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISOb_118.GSR = "DISABLED";
    LUT4 mux_9_i30_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[29]), .C(\speed_m4[17] ), 
         .D(n22202), .Z(MISOb_N_666[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 MISOb_N_667_bdd_2_lut (.A(MISO_N_624), .B(MISO_N_625), .Z(n21481)) /* synthesis lut_function=(A (B)) */ ;
    defparam MISOb_N_667_bdd_2_lut.init = 16'h8888;
    LUT4 mux_9_i31_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[30]), .C(\speed_m4[18] ), 
         .D(n22202), .Z(MISOb_N_666[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i13588_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[31]), .C(\speed_m4[19] ), 
         .D(n22202), .Z(MISOb_N_666[31])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam i13588_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i34_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[33]), .C(\speed_m3[0] ), 
         .D(n22202), .Z(MISOb_N_666[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i35_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[34]), .C(\speed_m3[1] ), 
         .D(n22202), .Z(MISOb_N_666[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i36_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[35]), .C(\speed_m3[2] ), 
         .D(n22202), .Z(MISOb_N_666[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i37_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[36]), .C(\speed_m3[3] ), 
         .D(n22202), .Z(MISOb_N_666[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i38_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[37]), .C(\speed_m3[4] ), 
         .D(n22202), .Z(MISOb_N_666[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX \SPI__7__i83  (.D(MOSI_c), .SP(clkout_c_enable_61), .CK(clkout_c), 
            .Q(recv_buffer[95]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i83 .GSR = "DISABLED";
    LUT4 mux_9_i39_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[38]), .C(\speed_m3[5] ), 
         .D(n22202), .Z(MISOb_N_666[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i40_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[39]), .C(\speed_m3[6] ), 
         .D(n22202), .Z(MISOb_N_666[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i41_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[40]), .C(\speed_m3[7] ), 
         .D(n22202), .Z(MISOb_N_666[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i10_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[9]), .C(enable_m3), 
         .D(n22202), .Z(MISOb_N_666[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i9_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[8]), .C(enable_m4), 
         .D(n22202), .Z(MISOb_N_666[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i42_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[41]), .C(\speed_m3[8] ), 
         .D(n22202), .Z(MISOb_N_666[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i43_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[42]), .C(\speed_m3[9] ), 
         .D(n22202), .Z(MISOb_N_666[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 MISOb_N_667_bdd_4_lut (.A(n21580), .B(send_buffer[1]), .C(MISOb), 
         .D(n21555), .Z(n21480)) /* synthesis lut_function=(A (B+(D))+!A !((D)+!C)) */ ;
    defparam MISOb_N_667_bdd_4_lut.init = 16'haad8;
    LUT4 mux_9_i44_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[43]), .C(\speed_m3[10] ), 
         .D(n22202), .Z(MISOb_N_666[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i45_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[44]), .C(\speed_m3[11] ), 
         .D(n22202), .Z(MISOb_N_666[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i46_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[45]), .C(\speed_m3[12] ), 
         .D(n22202), .Z(MISOb_N_666[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i47_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[46]), .C(\speed_m3[13] ), 
         .D(n22202), .Z(MISOb_N_666[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i48_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[47]), .C(\speed_m3[14] ), 
         .D(n22202), .Z(MISOb_N_666[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i49_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[48]), .C(\speed_m3[15] ), 
         .D(n22202), .Z(MISOb_N_666[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i50_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[49]), .C(\speed_m3[16] ), 
         .D(n22202), .Z(MISOb_N_666[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i51_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[50]), .C(\speed_m3[17] ), 
         .D(n22202), .Z(MISOb_N_666[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i52_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[51]), .C(\speed_m3[18] ), 
         .D(n22202), .Z(MISOb_N_666[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i13587_3_lut_4_lut_4_lut (.A(CSlatched), .B(send_buffer[52]), .C(\speed_m3[19] ), 
         .D(CSold), .Z(MISOb_N_666[52])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam i13587_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i55_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[54]), .C(\speed_m2[0] ), 
         .D(n22202), .Z(MISOb_N_666[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i56_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[55]), .C(\speed_m2[1] ), 
         .D(n22202), .Z(MISOb_N_666[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i57_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[56]), .C(\speed_m2[2] ), 
         .D(n22202), .Z(MISOb_N_666[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i58_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[57]), .C(\speed_m2[3] ), 
         .D(n22202), .Z(MISOb_N_666[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i59_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[58]), .C(\speed_m2[4] ), 
         .D(n22202), .Z(MISOb_N_666[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX \SPI__7__i82  (.D(recv_buffer[95]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[94]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i82 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i81  (.D(recv_buffer[94]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[93]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i81 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i80  (.D(recv_buffer[93]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[92]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i80 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i79  (.D(recv_buffer[92]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[91]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i79 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i78  (.D(recv_buffer[91]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[90]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i78 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i77  (.D(recv_buffer[90]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[89]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i77 .GSR = "DISABLED";
    LUT4 mux_9_i60_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[59]), .C(\speed_m2[5] ), 
         .D(n22202), .Z(MISOb_N_666[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i18_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[17]), .C(\speed_m4[5] ), 
         .D(n22202), .Z(MISOb_N_666[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX \SPI__7__i76  (.D(recv_buffer[89]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[88]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i76 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i75  (.D(recv_buffer[88]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[87]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i75 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i74  (.D(recv_buffer[87]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[86]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i74 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i73  (.D(recv_buffer[86]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[85]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i73 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i72  (.D(recv_buffer[85]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[84]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i72 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i71  (.D(recv_buffer[84]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[83]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i71 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i70  (.D(recv_buffer[83]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[82]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i70 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i69  (.D(recv_buffer[82]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[81]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i69 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i68  (.D(recv_buffer[81]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[80]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i68 .GSR = "DISABLED";
    LUT4 mux_9_i17_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[16]), .C(\speed_m4[4] ), 
         .D(n22202), .Z(MISOb_N_666[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i61_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[60]), .C(\speed_m2[6] ), 
         .D(n22202), .Z(MISOb_N_666[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i62_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[61]), .C(\speed_m2[7] ), 
         .D(n22202), .Z(MISOb_N_666[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i63_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[62]), .C(\speed_m2[8] ), 
         .D(n22202), .Z(MISOb_N_666[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i64_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[63]), .C(\speed_m2[9] ), 
         .D(n22202), .Z(MISOb_N_666[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i65_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[64]), .C(\speed_m2[10] ), 
         .D(n22202), .Z(MISOb_N_666[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i66_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[65]), .C(\speed_m2[11] ), 
         .D(n22202), .Z(MISOb_N_666[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i67_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[66]), .C(\speed_m2[12] ), 
         .D(n22202), .Z(MISOb_N_666[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i68_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[67]), .C(\speed_m2[13] ), 
         .D(n22202), .Z(MISOb_N_666[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i69_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[68]), .C(\speed_m2[14] ), 
         .D(n22202), .Z(MISOb_N_666[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i70_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[69]), .C(\speed_m2[15] ), 
         .D(n22202), .Z(MISOb_N_666[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i71_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[70]), .C(\speed_m2[16] ), 
         .D(n22202), .Z(MISOb_N_666[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i72_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[71]), .C(\speed_m2[17] ), 
         .D(n22202), .Z(MISOb_N_666[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i73_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[72]), .C(\speed_m2[18] ), 
         .D(n22202), .Z(MISOb_N_666[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i13586_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[73]), .C(\speed_m2[19] ), 
         .D(n22202), .Z(MISOb_N_666[73])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam i13586_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i76_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[75]), .C(\speed_m1[0] ), 
         .D(n22202), .Z(MISOb_N_666[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i77_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[76]), .C(\speed_m1[1] ), 
         .D(n22202), .Z(MISOb_N_666[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i78_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[77]), .C(\speed_m1[2] ), 
         .D(n22202), .Z(MISOb_N_666[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i79_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[78]), .C(\speed_m1[3] ), 
         .D(n22202), .Z(MISOb_N_666[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i80_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[79]), .C(\speed_m1[4] ), 
         .D(n22202), .Z(MISOb_N_666[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i20_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[19]), .C(\speed_m4[7] ), 
         .D(n22202), .Z(MISOb_N_666[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i19_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[18]), .C(\speed_m4[6] ), 
         .D(n22202), .Z(MISOb_N_666[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i81_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[80]), .C(\speed_m1[5] ), 
         .D(n22202), .Z(MISOb_N_666[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i82_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[81]), .C(\speed_m1[6] ), 
         .D(n22202), .Z(MISOb_N_666[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i83_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[82]), .C(\speed_m1[7] ), 
         .D(n22202), .Z(MISOb_N_666[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i84_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[83]), .C(\speed_m1[8] ), 
         .D(n22202), .Z(MISOb_N_666[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i85_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[84]), .C(\speed_m1[9] ), 
         .D(n22202), .Z(MISOb_N_666[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i86_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[85]), .C(\speed_m1[10] ), 
         .D(n22202), .Z(MISOb_N_666[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i87_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[86]), .C(\speed_m1[11] ), 
         .D(n22202), .Z(MISOb_N_666[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i88_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[87]), .C(\speed_m1[12] ), 
         .D(n22202), .Z(MISOb_N_666[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i89_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[88]), .C(\speed_m1[13] ), 
         .D(n22202), .Z(MISOb_N_666[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i90_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[89]), .C(\speed_m1[14] ), 
         .D(n22202), .Z(MISOb_N_666[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i91_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[90]), .C(\speed_m1[15] ), 
         .D(n22202), .Z(MISOb_N_666[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i92_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[91]), .C(\speed_m1[16] ), 
         .D(n22202), .Z(MISOb_N_666[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i93_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[92]), .C(\speed_m1[17] ), 
         .D(n22202), .Z(MISOb_N_666[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i94_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[93]), .C(\speed_m1[18] ), 
         .D(n22202), .Z(MISOb_N_666[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i21_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[20]), .C(\speed_m4[8] ), 
         .D(n22202), .Z(MISOb_N_666[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i11_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[10]), .C(enable_m2), 
         .D(n22202), .Z(MISOb_N_666[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i12_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[11]), .C(enable_m1), 
         .D(n22202), .Z(MISOb_N_666[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i13575_3_lut_rep_316_4_lut_4_lut (.A(CSlatched), .B(\send_buffer[94] ), 
         .C(\speed_m1[19] ), .D(CSold), .Z(n21525)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam i13575_3_lut_rep_316_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i13_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[12]), .C(\speed_m4[0] ), 
         .D(n22202), .Z(MISOb_N_666[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i14_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[13]), .C(\speed_m4[1] ), 
         .D(n22202), .Z(MISOb_N_666[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i15_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[14]), .C(\speed_m4[2] ), 
         .D(n22202), .Z(MISOb_N_666[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX \SPI__7__i67  (.D(recv_buffer[80]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[79]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i67 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i66  (.D(recv_buffer[79]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[78]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i66 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i65  (.D(recv_buffer[78]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[77]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i65 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i64  (.D(recv_buffer[77]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[76]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i64 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i63  (.D(recv_buffer[76]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[75]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i63 .GSR = "DISABLED";
    LUT4 mux_9_i16_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[15]), .C(\speed_m4[3] ), 
         .D(n22202), .Z(MISOb_N_666[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i9_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[8]), 
         .C(MISOb_N_666[9]), .D(n21580), .Z(send_buffer_95__N_346[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i10_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[9]), 
         .C(MISOb_N_666[10]), .D(n21580), .Z(send_buffer_95__N_346[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX \SPI__7__i62  (.D(recv_buffer[75]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[74]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i62 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i61  (.D(recv_buffer[74]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[73]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i61 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i60  (.D(recv_buffer[73]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[72]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i60 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i59  (.D(recv_buffer[72]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[71]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i59 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i58  (.D(recv_buffer[71]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[70]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i58 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i57  (.D(recv_buffer[70]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[69]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i57 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i56  (.D(recv_buffer[69]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[68]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i56 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i55  (.D(recv_buffer[68]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[67]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i55 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i54  (.D(recv_buffer[67]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[66]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i54 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i53  (.D(recv_buffer[66]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[65]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i53 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i52  (.D(recv_buffer[65]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[64]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i52 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i51  (.D(recv_buffer[64]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[63]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i51 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i50  (.D(recv_buffer[63]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[62]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i50 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i49  (.D(recv_buffer[62]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[61]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i49 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i48  (.D(recv_buffer[61]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[60]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i48 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i47  (.D(recv_buffer[60]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[59]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i47 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i46  (.D(recv_buffer[59]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[58]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i46 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i45  (.D(recv_buffer[58]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[57]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i45 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i44  (.D(recv_buffer[57]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[56]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i44 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i43  (.D(recv_buffer[56]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[55]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i43 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i42  (.D(recv_buffer[55]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[54]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i42 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i41  (.D(recv_buffer[54]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[53]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i41 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i40  (.D(recv_buffer[53]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[52]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i40 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i39  (.D(recv_buffer[52]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[51]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i39 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i38  (.D(recv_buffer[51]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[50]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i38 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i37  (.D(recv_buffer[50]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[49]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i37 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i36  (.D(recv_buffer[49]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[48]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i36 .GSR = "DISABLED";
    LUT4 mux_51_i11_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[10]), 
         .C(MISOb_N_666[11]), .D(n21580), .Z(send_buffer_95__N_346[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX \SPI__7__i35  (.D(recv_buffer[48]), .SP(clkout_c_enable_61), 
            .CK(clkout_c), .Q(recv_buffer[47]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i35 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i34  (.D(recv_buffer[47]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[46]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i34 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i33  (.D(recv_buffer[46]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[45]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i33 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i32  (.D(recv_buffer[45]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[44]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i32 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i31  (.D(recv_buffer[44]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[43]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i31 .GSR = "DISABLED";
    LUT4 mux_51_i12_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[11]), 
         .C(MISOb_N_666[12]), .D(n21580), .Z(send_buffer_95__N_346[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX \SPI__7__i30  (.D(recv_buffer[43]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[42]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i30 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i29  (.D(recv_buffer[42]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[41]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i29 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i28  (.D(recv_buffer[41]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[40]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i28 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i27  (.D(recv_buffer[40]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[39]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i27 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i26  (.D(recv_buffer[39]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[38]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i26 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i25  (.D(recv_buffer[38]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[37]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i25 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i24  (.D(recv_buffer[37]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[36]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i24 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i23  (.D(recv_buffer[36]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[35]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i23 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i22  (.D(recv_buffer[35]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[34]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i22 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i21  (.D(recv_buffer[34]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[33]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i21 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i20  (.D(recv_buffer[33]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[32]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i20 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i19  (.D(recv_buffer[32]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[31]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i19 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i18  (.D(recv_buffer[31]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[30]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i18 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i17  (.D(recv_buffer[30]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[29]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i17 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i16  (.D(recv_buffer[29]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[28]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i16 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i15  (.D(recv_buffer[28]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[27]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i15 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i14  (.D(recv_buffer[27]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[26]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i14 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i13  (.D(recv_buffer[26]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[25]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i13 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i12  (.D(recv_buffer[25]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[24]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i12 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i11  (.D(recv_buffer[24]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[23]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i11 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i10  (.D(recv_buffer[23]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[22]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i10 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i9  (.D(recv_buffer[22]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[21]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i9 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i8  (.D(recv_buffer[21]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[20]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i8 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i7  (.D(recv_buffer[20]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[19]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i7 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i6  (.D(recv_buffer[19]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i6 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i5  (.D(recv_buffer[18]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[17]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i5 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i4  (.D(recv_buffer[17]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i4 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i3  (.D(recv_buffer[16]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[15]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i3 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i2  (.D(recv_buffer[15]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i2 .GSR = "DISABLED";
    FD1P3AX \SPI__7__i1  (.D(recv_buffer[14]), .SP(clkout_c_enable_96), 
            .CK(clkout_c), .Q(recv_buffer[13]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__7__i1 .GSR = "DISABLED";
    LUT4 mux_51_i13_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[12]), 
         .C(MISOb_N_666[13]), .D(n21580), .Z(send_buffer_95__N_346[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i14_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[13]), 
         .C(MISOb_N_666[14]), .D(n21580), .Z(send_buffer_95__N_346[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i15_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[14]), 
         .C(MISOb_N_666[15]), .D(n21580), .Z(send_buffer_95__N_346[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i16_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[15]), 
         .C(MISOb_N_666[16]), .D(n21580), .Z(send_buffer_95__N_346[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i17_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[16]), 
         .C(MISOb_N_666[17]), .D(n21580), .Z(send_buffer_95__N_346[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i18_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[17]), 
         .C(MISOb_N_666[18]), .D(n21580), .Z(send_buffer_95__N_346[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i19_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[18]), 
         .C(MISOb_N_666[19]), .D(n21580), .Z(send_buffer_95__N_346[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i20_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[19]), 
         .C(MISOb_N_666[20]), .D(n21580), .Z(send_buffer_95__N_346[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i21_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[20]), 
         .C(MISOb_N_666[21]), .D(n21580), .Z(send_buffer_95__N_346[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i22_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[21]), 
         .C(MISOb_N_666[22]), .D(n21580), .Z(send_buffer_95__N_346[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i23_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[22]), 
         .C(MISOb_N_666[23]), .D(n21580), .Z(send_buffer_95__N_346[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i24_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[23]), 
         .C(MISOb_N_666[24]), .D(n21580), .Z(send_buffer_95__N_346[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i25_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[24]), 
         .C(MISOb_N_666[25]), .D(n21580), .Z(send_buffer_95__N_346[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i26_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[25]), 
         .C(MISOb_N_666[26]), .D(n21580), .Z(send_buffer_95__N_346[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3JX speed_set_m3_i0_i0 (.D(recv_buffer[33]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i0.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i0 (.D(recv_buffer[54]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i0.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i0 (.D(recv_buffer[75]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i0.GSR = "DISABLED";
    LUT4 mux_51_i27_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[26]), 
         .C(MISOb_N_666[27]), .D(n21580), .Z(send_buffer_95__N_346[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i28_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[27]), 
         .C(MISOb_N_666[28]), .D(n21580), .Z(send_buffer_95__N_346[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i29_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[28]), 
         .C(MISOb_N_666[29]), .D(n21580), .Z(send_buffer_95__N_346[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i30_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[29]), 
         .C(MISOb_N_666[30]), .D(n21580), .Z(send_buffer_95__N_346[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i31_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[30]), 
         .C(MISOb_N_666[31]), .D(n21580), .Z(send_buffer_95__N_346[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i34_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[33]), 
         .C(MISOb_N_666[34]), .D(n21580), .Z(send_buffer_95__N_346[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i35_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[34]), 
         .C(MISOb_N_666[35]), .D(n21580), .Z(send_buffer_95__N_346[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i36_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[35]), 
         .C(MISOb_N_666[36]), .D(n21580), .Z(send_buffer_95__N_346[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i37_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[36]), 
         .C(MISOb_N_666[37]), .D(n21580), .Z(send_buffer_95__N_346[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i38_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[37]), 
         .C(MISOb_N_666[38]), .D(n21580), .Z(send_buffer_95__N_346[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i39_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[38]), 
         .C(MISOb_N_666[39]), .D(n21580), .Z(send_buffer_95__N_346[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i40_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[39]), 
         .C(MISOb_N_666[40]), .D(n21580), .Z(send_buffer_95__N_346[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i41_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[40]), 
         .C(MISOb_N_666[41]), .D(n21580), .Z(send_buffer_95__N_346[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i42_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[41]), 
         .C(MISOb_N_666[42]), .D(n21580), .Z(send_buffer_95__N_346[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i43_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[42]), 
         .C(MISOb_N_666[43]), .D(n21580), .Z(send_buffer_95__N_346[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i44_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[43]), 
         .C(MISOb_N_666[44]), .D(n21580), .Z(send_buffer_95__N_346[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i45_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[44]), 
         .C(MISOb_N_666[45]), .D(n21580), .Z(send_buffer_95__N_346[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i46_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[45]), 
         .C(MISOb_N_666[46]), .D(n21580), .Z(send_buffer_95__N_346[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i47_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[46]), 
         .C(MISOb_N_666[47]), .D(n21580), .Z(send_buffer_95__N_346[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i48_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[47]), 
         .C(MISOb_N_666[48]), .D(n21580), .Z(send_buffer_95__N_346[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i49_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[48]), 
         .C(MISOb_N_666[49]), .D(n21580), .Z(send_buffer_95__N_346[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i50_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[49]), 
         .C(MISOb_N_666[50]), .D(n21580), .Z(send_buffer_95__N_346[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 CSold_I_0_132_2_lut (.A(CSold), .B(CSlatched), .Z(enable_m1_N_633)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(139[7:42])
    defparam CSold_I_0_132_2_lut.init = 16'h8888;
    LUT4 mux_51_i51_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[50]), 
         .C(MISOb_N_666[51]), .D(n21580), .Z(send_buffer_95__N_346[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i52_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[51]), 
         .C(MISOb_N_666[52]), .D(n21580), .Z(send_buffer_95__N_346[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i55_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[54]), 
         .C(MISOb_N_666[55]), .D(n21580), .Z(send_buffer_95__N_346[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i56_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[55]), 
         .C(MISOb_N_666[56]), .D(n21580), .Z(send_buffer_95__N_346[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i57_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[56]), 
         .C(MISOb_N_666[57]), .D(n21580), .Z(send_buffer_95__N_346[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i58_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[57]), 
         .C(MISOb_N_666[58]), .D(n21580), .Z(send_buffer_95__N_346[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i59_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[58]), 
         .C(MISOb_N_666[59]), .D(n21580), .Z(send_buffer_95__N_346[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i60_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[59]), 
         .C(MISOb_N_666[60]), .D(n21580), .Z(send_buffer_95__N_346[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i61_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[60]), 
         .C(MISOb_N_666[61]), .D(n21580), .Z(send_buffer_95__N_346[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i62_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[61]), 
         .C(MISOb_N_666[62]), .D(n21580), .Z(send_buffer_95__N_346[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i63_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[62]), 
         .C(MISOb_N_666[63]), .D(n21580), .Z(send_buffer_95__N_346[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i64_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[63]), 
         .C(MISOb_N_666[64]), .D(n21580), .Z(send_buffer_95__N_346[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i2_4_lut (.A(n3479), .B(n3455), .C(n39_adj_1886), .D(n40_adj_1887), 
         .Z(enable_m4_N_649)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i18_4_lut (.A(recv_buffer[25]), .B(n36_adj_1888), .C(n28_adj_1889), 
         .D(recv_buffer[24]), .Z(n39_adj_1886)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 mux_51_i65_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[64]), 
         .C(MISOb_N_666[65]), .D(n21580), .Z(send_buffer_95__N_346[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i66_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[65]), 
         .C(MISOb_N_666[66]), .D(n21580), .Z(send_buffer_95__N_346[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i67_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[66]), 
         .C(MISOb_N_666[67]), .D(n21580), .Z(send_buffer_95__N_346[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i19_4_lut (.A(recv_buffer[27]), .B(n38_adj_1890), .C(n32_adj_1891), 
         .D(recv_buffer[22]), .Z(n40_adj_1887)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(n169[0]), .B(recv_buffer[19]), .C(recv_buffer[29]), 
         .D(recv_buffer[23]), .Z(n36_adj_1888)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 mux_51_i68_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[67]), 
         .C(MISOb_N_666[68]), .D(n21580), .Z(send_buffer_95__N_346[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i69_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[68]), 
         .C(MISOb_N_666[69]), .D(n21580), .Z(send_buffer_95__N_346[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i70_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[69]), 
         .C(MISOb_N_666[70]), .D(n21580), .Z(send_buffer_95__N_346[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i71_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[70]), 
         .C(MISOb_N_666[71]), .D(n21580), .Z(send_buffer_95__N_346[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i72_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[71]), 
         .C(MISOb_N_666[72]), .D(n21580), .Z(send_buffer_95__N_346[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i73_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[72]), 
         .C(MISOb_N_666[73]), .D(n21580), .Z(send_buffer_95__N_346[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i76_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[75]), 
         .C(MISOb_N_666[76]), .D(n21580), .Z(send_buffer_95__N_346[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i77_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[76]), 
         .C(MISOb_N_666[77]), .D(n21580), .Z(send_buffer_95__N_346[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i78_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[77]), 
         .C(MISOb_N_666[78]), .D(n21580), .Z(send_buffer_95__N_346[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i79_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[78]), 
         .C(MISOb_N_666[79]), .D(n21580), .Z(send_buffer_95__N_346[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i80_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[79]), 
         .C(MISOb_N_666[80]), .D(n21580), .Z(send_buffer_95__N_346[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i81_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[80]), 
         .C(MISOb_N_666[81]), .D(n21580), .Z(send_buffer_95__N_346[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i82_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[81]), 
         .C(MISOb_N_666[82]), .D(n21580), .Z(send_buffer_95__N_346[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i83_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[82]), 
         .C(MISOb_N_666[83]), .D(n21580), .Z(send_buffer_95__N_346[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i84_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[83]), 
         .C(MISOb_N_666[84]), .D(n21580), .Z(send_buffer_95__N_346[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i85_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[84]), 
         .C(MISOb_N_666[85]), .D(n21580), .Z(send_buffer_95__N_346[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i86_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[85]), 
         .C(MISOb_N_666[86]), .D(n21580), .Z(send_buffer_95__N_346[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i87_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[86]), 
         .C(MISOb_N_666[87]), .D(n21580), .Z(send_buffer_95__N_346[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i88_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[87]), 
         .C(MISOb_N_666[88]), .D(n21580), .Z(send_buffer_95__N_346[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i89_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[88]), 
         .C(MISOb_N_666[89]), .D(n21580), .Z(send_buffer_95__N_346[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i90_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[89]), 
         .C(MISOb_N_666[90]), .D(n21580), .Z(send_buffer_95__N_346[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i91_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[90]), 
         .C(MISOb_N_666[91]), .D(n21580), .Z(send_buffer_95__N_346[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i92_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[91]), 
         .C(MISOb_N_666[92]), .D(n21580), .Z(send_buffer_95__N_346[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i93_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[92]), 
         .C(MISOb_N_666[93]), .D(n21580), .Z(send_buffer_95__N_346[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i94_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_666[93]), 
         .C(n21525), .D(n21580), .Z(send_buffer_95__N_346[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_51_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i1_2_lut_rep_379 (.A(enable_m4), .B(free_m4), .Z(n21588)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_379.init = 16'h2222;
    LUT4 i17955_3_lut_4_lut (.A(enable_m4), .B(free_m4), .C(hallsense_m4[2]), 
         .D(hallsense_m4[0]), .Z(n19662)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17955_3_lut_4_lut.init = 16'hfddf;
    LUT4 i7_2_lut (.A(recv_buffer[13]), .B(recv_buffer[14]), .Z(n28_adj_1889)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_rep_410 (.A(SCKold), .B(n22203), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_61)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut_rep_410.init = 16'h0400;
    LUT4 mux_9_i25_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[24]), .C(\speed_m4[12] ), 
         .D(n22202), .Z(MISOb_N_666[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i17_4_lut (.A(recv_buffer[20]), .B(n34_adj_1892), .C(n24_adj_1893), 
         .D(recv_buffer[28]), .Z(n38_adj_1890)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    CCU2D add_15805_16 (.A0(recv_buffer[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18634), .S1(n3431));
    defparam add_15805_16.INIT0 = 16'h0aaa;
    defparam add_15805_16.INIT1 = 16'h0000;
    defparam add_15805_16.INJECT1_0 = "NO";
    defparam add_15805_16.INJECT1_1 = "NO";
    CCU2D add_15805_14 (.A0(recv_buffer[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18633), .COUT(n18634));
    defparam add_15805_14.INIT0 = 16'h5aaa;
    defparam add_15805_14.INIT1 = 16'h5aaa;
    defparam add_15805_14.INJECT1_0 = "NO";
    defparam add_15805_14.INJECT1_1 = "NO";
    CCU2D add_15805_12 (.A0(recv_buffer[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18632), .COUT(n18633));
    defparam add_15805_12.INIT0 = 16'h5aaa;
    defparam add_15805_12.INIT1 = 16'h5aaa;
    defparam add_15805_12.INJECT1_0 = "NO";
    defparam add_15805_12.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(recv_buffer[18]), .B(recv_buffer[15]), .C(recv_buffer[26]), 
         .Z(n32_adj_1891)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(recv_buffer[32]), .B(recv_buffer[31]), .C(recv_buffer[21]), 
         .D(recv_buffer[16]), .Z(n34_adj_1892)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(recv_buffer[30]), .B(recv_buffer[17]), .Z(n24_adj_1893)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    FD1P3AX send_buffer_i0_i1 (.D(send_buffer_95__N_346[1]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i1.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i2 (.D(send_buffer_95__N_346[2]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i3 (.D(send_buffer_95__N_346[3]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i4 (.D(send_buffer_95__N_346[4]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i4.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i5 (.D(send_buffer_95__N_346[5]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i5.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i6 (.D(send_buffer_95__N_346[6]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i7 (.D(send_buffer_95__N_346[7]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i8 (.D(send_buffer_95__N_346[8]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i8.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i9 (.D(send_buffer_95__N_346[9]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i9.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i10 (.D(send_buffer_95__N_346[10]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i10.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i11 (.D(send_buffer_95__N_346[11]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i11.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i12 (.D(send_buffer_95__N_346[12]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i12.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i13 (.D(send_buffer_95__N_346[13]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i13.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i14 (.D(send_buffer_95__N_346[14]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i14.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i15 (.D(send_buffer_95__N_346[15]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i15.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i16 (.D(send_buffer_95__N_346[16]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i16.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i17 (.D(send_buffer_95__N_346[17]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i17.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i18 (.D(send_buffer_95__N_346[18]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i18.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i19 (.D(send_buffer_95__N_346[19]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i19.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i20 (.D(send_buffer_95__N_346[20]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i20.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i21 (.D(send_buffer_95__N_346[21]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i21.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i22 (.D(send_buffer_95__N_346[22]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i22.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i23 (.D(send_buffer_95__N_346[23]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i23.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i24 (.D(send_buffer_95__N_346[24]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i24.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i25 (.D(send_buffer_95__N_346[25]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i25.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i26 (.D(send_buffer_95__N_346[26]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i26.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i27 (.D(send_buffer_95__N_346[27]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i27.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i28 (.D(send_buffer_95__N_346[28]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i28.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i29 (.D(send_buffer_95__N_346[29]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i29.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i30 (.D(send_buffer_95__N_346[30]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i30.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i31 (.D(send_buffer_95__N_346[31]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i31.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i32 (.D(send_buffer_95__N_346[32]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i32.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i33 (.D(send_buffer_95__N_346[33]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i33.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i34 (.D(send_buffer_95__N_346[34]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i34.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i35 (.D(send_buffer_95__N_346[35]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i35.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i36 (.D(send_buffer_95__N_346[36]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i36.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i37 (.D(send_buffer_95__N_346[37]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i37.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i38 (.D(send_buffer_95__N_346[38]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i38.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i39 (.D(send_buffer_95__N_346[39]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i39.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i40 (.D(send_buffer_95__N_346[40]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i40.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i41 (.D(send_buffer_95__N_346[41]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i41.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i42 (.D(send_buffer_95__N_346[42]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i42.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i43 (.D(send_buffer_95__N_346[43]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i43.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i44 (.D(send_buffer_95__N_346[44]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i44.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i45 (.D(send_buffer_95__N_346[45]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i45.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i46 (.D(send_buffer_95__N_346[46]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i46.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i47 (.D(send_buffer_95__N_346[47]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i47.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i48 (.D(send_buffer_95__N_346[48]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i48.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i49 (.D(send_buffer_95__N_346[49]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i49.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i50 (.D(send_buffer_95__N_346[50]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i50.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i51 (.D(send_buffer_95__N_346[51]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i51.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i52 (.D(send_buffer_95__N_346[52]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i52.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i53 (.D(send_buffer_95__N_346[53]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i53.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i54 (.D(send_buffer_95__N_346[54]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i54.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i55 (.D(send_buffer_95__N_346[55]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i55.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i56 (.D(send_buffer_95__N_346[56]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i56.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i57 (.D(send_buffer_95__N_346[57]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i57.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i58 (.D(send_buffer_95__N_346[58]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i58.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i59 (.D(send_buffer_95__N_346[59]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i59.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i60 (.D(send_buffer_95__N_346[60]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i60.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i61 (.D(send_buffer_95__N_346[61]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i61.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i62 (.D(send_buffer_95__N_346[62]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i62.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i63 (.D(send_buffer_95__N_346[63]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i63.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i64 (.D(send_buffer_95__N_346[64]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i64.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i65 (.D(send_buffer_95__N_346[65]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i65.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i66 (.D(send_buffer_95__N_346[66]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i66.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i67 (.D(send_buffer_95__N_346[67]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i67.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i68 (.D(send_buffer_95__N_346[68]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i68.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i69 (.D(send_buffer_95__N_346[69]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i69.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i70 (.D(send_buffer_95__N_346[70]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i70.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i71 (.D(send_buffer_95__N_346[71]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i71.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i72 (.D(send_buffer_95__N_346[72]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i72.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i73 (.D(send_buffer_95__N_346[73]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i73.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i74 (.D(send_buffer_95__N_346[74]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i74.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i75 (.D(send_buffer_95__N_346[75]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i75.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i76 (.D(send_buffer_95__N_346[76]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i76.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i77 (.D(send_buffer_95__N_346[77]), .SP(clkout_c_enable_176), 
            .CK(clkout_c), .Q(send_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i77.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i78 (.D(send_buffer_95__N_346[78]), .SP(clkout_c_enable_164), 
            .CK(clkout_c), .Q(send_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i78.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i79 (.D(send_buffer_95__N_346[79]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i79.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i80 (.D(send_buffer_95__N_346[80]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i80.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i81 (.D(send_buffer_95__N_346[81]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i81.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i82 (.D(send_buffer_95__N_346[82]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i82.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i83 (.D(send_buffer_95__N_346[83]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i83.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i84 (.D(send_buffer_95__N_346[84]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i84.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i85 (.D(send_buffer_95__N_346[85]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i85.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i86 (.D(send_buffer_95__N_346[86]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i86.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i87 (.D(send_buffer_95__N_346[87]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i87.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i88 (.D(send_buffer_95__N_346[88]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i88.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i89 (.D(send_buffer_95__N_346[89]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i89.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i90 (.D(send_buffer_95__N_346[90]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i90.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i91 (.D(send_buffer_95__N_346[91]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i91.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i92 (.D(send_buffer_95__N_346[92]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i92.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i93 (.D(send_buffer_95__N_346[93]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i93.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i94 (.D(\send_buffer_95__N_346[94] ), .SP(rst), 
            .CK(clkout_c), .Q(\send_buffer[94] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i94.GSR = "DISABLED";
    CCU2D add_15805_10 (.A0(recv_buffer[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18631), .COUT(n18632));
    defparam add_15805_10.INIT0 = 16'h5555;
    defparam add_15805_10.INIT1 = 16'h5aaa;
    defparam add_15805_10.INJECT1_0 = "NO";
    defparam add_15805_10.INJECT1_1 = "NO";
    CCU2D add_15805_8 (.A0(recv_buffer[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18630), .COUT(n18631));
    defparam add_15805_8.INIT0 = 16'h5aaa;
    defparam add_15805_8.INIT1 = 16'h5aaa;
    defparam add_15805_8.INJECT1_0 = "NO";
    defparam add_15805_8.INJECT1_1 = "NO";
    CCU2D add_15805_6 (.A0(recv_buffer[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18629), .COUT(n18630));
    defparam add_15805_6.INIT0 = 16'h5555;
    defparam add_15805_6.INIT1 = 16'h5555;
    defparam add_15805_6.INJECT1_0 = "NO";
    defparam add_15805_6.INJECT1_1 = "NO";
    CCU2D add_15805_4 (.A0(recv_buffer[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18628), .COUT(n18629));
    defparam add_15805_4.INIT0 = 16'h5aaa;
    defparam add_15805_4.INIT1 = 16'h5555;
    defparam add_15805_4.INJECT1_0 = "NO";
    defparam add_15805_4.INJECT1_1 = "NO";
    CCU2D add_15805_2 (.A0(recv_buffer[39]), .B0(recv_buffer[38]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18628));
    defparam add_15805_2.INIT0 = 16'h7000;
    defparam add_15805_2.INIT1 = 16'h5aaa;
    defparam add_15805_2.INJECT1_0 = "NO";
    defparam add_15805_2.INJECT1_1 = "NO";
    CCU2D add_15806_16 (.A0(recv_buffer[74]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18627), .S1(n3383));
    defparam add_15806_16.INIT0 = 16'h0aaa;
    defparam add_15806_16.INIT1 = 16'h0000;
    defparam add_15806_16.INJECT1_0 = "NO";
    defparam add_15806_16.INJECT1_1 = "NO";
    CCU2D add_15806_14 (.A0(recv_buffer[72]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[73]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18626), .COUT(n18627));
    defparam add_15806_14.INIT0 = 16'h5aaa;
    defparam add_15806_14.INIT1 = 16'h5aaa;
    defparam add_15806_14.INJECT1_0 = "NO";
    defparam add_15806_14.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_388 (.A(enable_m2), .B(free_m2), .Z(n21597)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_388.init = 16'h2222;
    CCU2D add_15806_12 (.A0(recv_buffer[70]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[71]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18625), .COUT(n18626));
    defparam add_15806_12.INIT0 = 16'h5aaa;
    defparam add_15806_12.INIT1 = 16'h5aaa;
    defparam add_15806_12.INJECT1_0 = "NO";
    defparam add_15806_12.INJECT1_1 = "NO";
    CCU2D add_15806_10 (.A0(recv_buffer[68]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[69]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18624), .COUT(n18625));
    defparam add_15806_10.INIT0 = 16'h5555;
    defparam add_15806_10.INIT1 = 16'h5aaa;
    defparam add_15806_10.INJECT1_0 = "NO";
    defparam add_15806_10.INJECT1_1 = "NO";
    CCU2D add_15806_8 (.A0(recv_buffer[66]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[67]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18623), .COUT(n18624));
    defparam add_15806_8.INIT0 = 16'h5aaa;
    defparam add_15806_8.INIT1 = 16'h5aaa;
    defparam add_15806_8.INJECT1_0 = "NO";
    defparam add_15806_8.INJECT1_1 = "NO";
    LUT4 i17935_3_lut_4_lut (.A(enable_m2), .B(free_m2), .C(hallsense_m2[2]), 
         .D(hallsense_m2[0]), .Z(n19656)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17935_3_lut_4_lut.init = 16'hfddf;
    CCU2D add_15806_6 (.A0(recv_buffer[64]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[65]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18622), .COUT(n18623));
    defparam add_15806_6.INIT0 = 16'h5555;
    defparam add_15806_6.INIT1 = 16'h5555;
    defparam add_15806_6.INJECT1_0 = "NO";
    defparam add_15806_6.INJECT1_1 = "NO";
    CCU2D add_15806_4 (.A0(recv_buffer[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18621), .COUT(n18622));
    defparam add_15806_4.INIT0 = 16'h5aaa;
    defparam add_15806_4.INIT1 = 16'h5555;
    defparam add_15806_4.INJECT1_0 = "NO";
    defparam add_15806_4.INJECT1_1 = "NO";
    LUT4 i2655_1_lut (.A(MISO_N_625), .Z(n4883)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(64[1] 216[13])
    defparam i2655_1_lut.init = 16'h5555;
    CCU2D add_15806_2 (.A0(recv_buffer[60]), .B0(recv_buffer[59]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18621));
    defparam add_15806_2.INIT0 = 16'h7000;
    defparam add_15806_2.INIT1 = 16'h5aaa;
    defparam add_15806_2.INJECT1_0 = "NO";
    defparam add_15806_2.INJECT1_1 = "NO";
    CCU2D add_15807_21 (.A0(recv_buffer[74]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18620), .S1(n3359));
    defparam add_15807_21.INIT0 = 16'h5555;
    defparam add_15807_21.INIT1 = 16'h0000;
    defparam add_15807_21.INJECT1_0 = "NO";
    defparam add_15807_21.INJECT1_1 = "NO";
    CCU2D add_15807_19 (.A0(recv_buffer[72]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[73]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18619), .COUT(n18620));
    defparam add_15807_19.INIT0 = 16'hf555;
    defparam add_15807_19.INIT1 = 16'hf555;
    defparam add_15807_19.INJECT1_0 = "NO";
    defparam add_15807_19.INJECT1_1 = "NO";
    CCU2D add_15807_17 (.A0(recv_buffer[70]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[71]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18618), .COUT(n18619));
    defparam add_15807_17.INIT0 = 16'hf555;
    defparam add_15807_17.INIT1 = 16'hf555;
    defparam add_15807_17.INJECT1_0 = "NO";
    defparam add_15807_17.INJECT1_1 = "NO";
    CCU2D add_15807_15 (.A0(recv_buffer[68]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[69]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18617), .COUT(n18618));
    defparam add_15807_15.INIT0 = 16'h0aaa;
    defparam add_15807_15.INIT1 = 16'hf555;
    defparam add_15807_15.INJECT1_0 = "NO";
    defparam add_15807_15.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_395 (.A(CSlatched), .B(CSold), .C(n22203), .Z(clkout_c_enable_245)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(139[7:42])
    defparam i2_3_lut_rep_395.init = 16'h8080;
    LUT4 i10330_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22203), .D(enable_m1_N_627), 
         .Z(n12617)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(139[7:42])
    defparam i10330_2_lut_4_lut.init = 16'h0080;
    LUT4 i10310_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22203), .D(enable_m2_N_635), 
         .Z(n12597)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(139[7:42])
    defparam i10310_2_lut_4_lut.init = 16'h0080;
    LUT4 i10290_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22203), .D(enable_m3_N_642), 
         .Z(n12577)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(139[7:42])
    defparam i10290_2_lut_4_lut.init = 16'h0080;
    LUT4 i10270_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22203), .D(enable_m4_N_649), 
         .Z(n12557)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(139[7:42])
    defparam i10270_2_lut_4_lut.init = 16'h0080;
    CCU2D add_15807_13 (.A0(recv_buffer[66]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[67]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18616), .COUT(n18617));
    defparam add_15807_13.INIT0 = 16'hf555;
    defparam add_15807_13.INIT1 = 16'hf555;
    defparam add_15807_13.INJECT1_0 = "NO";
    defparam add_15807_13.INJECT1_1 = "NO";
    CCU2D add_15807_11 (.A0(recv_buffer[64]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[65]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18615), .COUT(n18616));
    defparam add_15807_11.INIT0 = 16'h0aaa;
    defparam add_15807_11.INIT1 = 16'h0aaa;
    defparam add_15807_11.INJECT1_0 = "NO";
    defparam add_15807_11.INJECT1_1 = "NO";
    CCU2D add_15807_9 (.A0(recv_buffer[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18614), .COUT(n18615));
    defparam add_15807_9.INIT0 = 16'hf555;
    defparam add_15807_9.INIT1 = 16'h0aaa;
    defparam add_15807_9.INJECT1_0 = "NO";
    defparam add_15807_9.INJECT1_1 = "NO";
    CCU2D add_15807_7 (.A0(recv_buffer[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18613), .COUT(n18614));
    defparam add_15807_7.INIT0 = 16'hf555;
    defparam add_15807_7.INIT1 = 16'hf555;
    defparam add_15807_7.INJECT1_0 = "NO";
    defparam add_15807_7.INJECT1_1 = "NO";
    CCU2D add_15807_5 (.A0(recv_buffer[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18612), .COUT(n18613));
    defparam add_15807_5.INIT0 = 16'hf555;
    defparam add_15807_5.INIT1 = 16'h0aaa;
    defparam add_15807_5.INJECT1_0 = "NO";
    defparam add_15807_5.INJECT1_1 = "NO";
    CCU2D add_15807_3 (.A0(recv_buffer[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18611), .COUT(n18612));
    defparam add_15807_3.INIT0 = 16'hf555;
    defparam add_15807_3.INIT1 = 16'hf555;
    defparam add_15807_3.INJECT1_0 = "NO";
    defparam add_15807_3.INJECT1_1 = "NO";
    CCU2D add_15807_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[54]), .B1(recv_buffer[55]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18611));
    defparam add_15807_1.INIT0 = 16'hF000;
    defparam add_15807_1.INIT1 = 16'ha666;
    defparam add_15807_1.INJECT1_0 = "NO";
    defparam add_15807_1.INJECT1_1 = "NO";
    CCU2D add_15808_16 (.A0(recv_buffer[95]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18610), .S1(n3335));
    defparam add_15808_16.INIT0 = 16'h0aaa;
    defparam add_15808_16.INIT1 = 16'h0000;
    defparam add_15808_16.INJECT1_0 = "NO";
    defparam add_15808_16.INJECT1_1 = "NO";
    CCU2D add_15808_14 (.A0(recv_buffer[93]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[94]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18609), .COUT(n18610));
    defparam add_15808_14.INIT0 = 16'h5aaa;
    defparam add_15808_14.INIT1 = 16'h5aaa;
    defparam add_15808_14.INJECT1_0 = "NO";
    defparam add_15808_14.INJECT1_1 = "NO";
    CCU2D add_15808_12 (.A0(recv_buffer[91]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[92]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18608), .COUT(n18609));
    defparam add_15808_12.INIT0 = 16'h5aaa;
    defparam add_15808_12.INIT1 = 16'h5aaa;
    defparam add_15808_12.INJECT1_0 = "NO";
    defparam add_15808_12.INJECT1_1 = "NO";
    CCU2D add_15808_10 (.A0(recv_buffer[89]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[90]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18607), .COUT(n18608));
    defparam add_15808_10.INIT0 = 16'h5555;
    defparam add_15808_10.INIT1 = 16'h5aaa;
    defparam add_15808_10.INJECT1_0 = "NO";
    defparam add_15808_10.INJECT1_1 = "NO";
    CCU2D add_15808_8 (.A0(recv_buffer[87]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[88]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18606), .COUT(n18607));
    defparam add_15808_8.INIT0 = 16'h5aaa;
    defparam add_15808_8.INIT1 = 16'h5aaa;
    defparam add_15808_8.INJECT1_0 = "NO";
    defparam add_15808_8.INJECT1_1 = "NO";
    FD1P3AX CSold_113_rep_405 (.D(n22201), .SP(clkout_c_enable_164), .CK(clkout_c), 
            .Q(n22202));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_113_rep_405.GSR = "DISABLED";
    CCU2D add_15808_6 (.A0(recv_buffer[85]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[86]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18605), .COUT(n18606));
    defparam add_15808_6.INIT0 = 16'h5555;
    defparam add_15808_6.INIT1 = 16'h5555;
    defparam add_15808_6.INJECT1_0 = "NO";
    defparam add_15808_6.INJECT1_1 = "NO";
    FD1P3JX speed_set_m1_i0_i1 (.D(recv_buffer[76]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i1.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i2 (.D(recv_buffer[77]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i2.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i3 (.D(recv_buffer[78]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i4 (.D(recv_buffer[79]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i4.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i5 (.D(recv_buffer[80]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i6 (.D(recv_buffer[81]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i7 (.D(recv_buffer[82]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i8 (.D(recv_buffer[83]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i9 (.D(recv_buffer[84]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i9.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i10 (.D(recv_buffer[85]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i11 (.D(recv_buffer[86]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i11.GSR = "DISABLED";
    LUT4 i2892_3_lut_4_lut_4_lut (.A(MISOb), .B(n21555), .C(n21556), .D(send_buffer[1]), 
         .Z(MISOb_N_660)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam i2892_3_lut_4_lut_4_lut.init = 16'hf2c2;
    LUT4 mux_51_i74_3_lut_4_lut (.A(send_buffer[74]), .B(n21555), .C(n21556), 
         .D(MISOb_N_666[73]), .Z(send_buffer_95__N_346[73])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i74_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_51_i75_3_lut_4_lut (.A(send_buffer[74]), .B(n21555), .C(n21556), 
         .D(MISOb_N_666[75]), .Z(send_buffer_95__N_346[74])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i75_3_lut_4_lut.init = 16'hf202;
    LUT4 mux_51_i53_3_lut_4_lut (.A(send_buffer[53]), .B(n21555), .C(n21556), 
         .D(MISOb_N_666[52]), .Z(send_buffer_95__N_346[52])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i53_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_51_i54_3_lut_4_lut (.A(send_buffer[53]), .B(n21555), .C(n21556), 
         .D(MISOb_N_666[54]), .Z(send_buffer_95__N_346[53])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i54_3_lut_4_lut.init = 16'hf202;
    LUT4 mux_9_i29_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[28]), .C(\speed_m4[16] ), 
         .D(n22202), .Z(MISOb_N_666[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_51_i32_3_lut_4_lut (.A(send_buffer[32]), .B(n21555), .C(n21556), 
         .D(MISOb_N_666[31]), .Z(send_buffer_95__N_346[31])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i32_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_51_i33_3_lut_4_lut (.A(send_buffer[32]), .B(n21555), .C(n21556), 
         .D(MISOb_N_666[33]), .Z(send_buffer_95__N_346[32])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i33_3_lut_4_lut.init = 16'hf202;
    LUT4 mux_51_i8_3_lut_4_lut (.A(send_buffer[7]), .B(n21555), .C(n21556), 
         .D(MISOb_N_666[8]), .Z(send_buffer_95__N_346[7])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i8_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_51_i7_3_lut_4_lut_4_lut (.A(send_buffer[6]), .B(n21555), .C(n21556), 
         .D(send_buffer[7]), .Z(send_buffer_95__N_346[6])) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i7_3_lut_4_lut_4_lut.init = 16'hf2c2;
    LUT4 mux_51_i6_3_lut_4_lut_4_lut (.A(send_buffer[5]), .B(n21555), .C(n21556), 
         .D(send_buffer[6]), .Z(send_buffer_95__N_346[5])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i6_3_lut_4_lut_4_lut.init = 16'h3e0e;
    LUT4 mux_51_i5_3_lut_4_lut_4_lut (.A(send_buffer[4]), .B(n21555), .C(n21556), 
         .D(send_buffer[5]), .Z(send_buffer_95__N_346[4])) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i5_3_lut_4_lut_4_lut.init = 16'hf2c2;
    LUT4 mux_51_i4_3_lut_4_lut_4_lut (.A(send_buffer[3]), .B(n21555), .C(n21556), 
         .D(send_buffer[4]), .Z(send_buffer_95__N_346[3])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i4_3_lut_4_lut_4_lut.init = 16'h3e0e;
    LUT4 mux_51_i2_3_lut_4_lut_4_lut (.A(send_buffer[2]), .B(n21555), .C(n21556), 
         .D(send_buffer[1]), .Z(send_buffer_95__N_346[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A (B (C)+!B (C+!(D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i2_3_lut_4_lut_4_lut.init = 16'h2f2c;
    LUT4 mux_51_i3_3_lut_4_lut_4_lut (.A(send_buffer[2]), .B(n21555), .C(n21556), 
         .D(send_buffer[3]), .Z(send_buffer_95__N_346[2])) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam mux_51_i3_3_lut_4_lut_4_lut.init = 16'hf2c2;
    CCU2D add_15808_4 (.A0(recv_buffer[83]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[84]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18604), .COUT(n18605));
    defparam add_15808_4.INIT0 = 16'h5aaa;
    defparam add_15808_4.INIT1 = 16'h5555;
    defparam add_15808_4.INJECT1_0 = "NO";
    defparam add_15808_4.INJECT1_1 = "NO";
    CCU2D add_15808_2 (.A0(recv_buffer[81]), .B0(recv_buffer[80]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[82]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18604));
    defparam add_15808_2.INIT0 = 16'h7000;
    defparam add_15808_2.INIT1 = 16'h5aaa;
    defparam add_15808_2.INJECT1_0 = "NO";
    defparam add_15808_2.INJECT1_1 = "NO";
    FD1P3AX CSlatched_115_rep_404 (.D(CS_c), .SP(clkout_c_enable_176), .CK(clkout_c), 
            .Q(n22201));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_115_rep_404.GSR = "DISABLED";
    CCU2D add_15809_21 (.A0(recv_buffer[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18603), .S1(n3407));
    defparam add_15809_21.INIT0 = 16'h5555;
    defparam add_15809_21.INIT1 = 16'h0000;
    defparam add_15809_21.INJECT1_0 = "NO";
    defparam add_15809_21.INJECT1_1 = "NO";
    FD1P3IX speed_set_m1_i0_i12 (.D(recv_buffer[87]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i12.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i13 (.D(recv_buffer[88]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i13.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i14 (.D(recv_buffer[89]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i15 (.D(recv_buffer[90]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i15.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i16 (.D(recv_buffer[91]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i16.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i17 (.D(recv_buffer[92]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i17.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i18 (.D(recv_buffer[93]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i18.GSR = "DISABLED";
    CCU2D add_15809_19 (.A0(recv_buffer[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18602), .COUT(n18603));
    defparam add_15809_19.INIT0 = 16'hf555;
    defparam add_15809_19.INIT1 = 16'hf555;
    defparam add_15809_19.INJECT1_0 = "NO";
    defparam add_15809_19.INJECT1_1 = "NO";
    CCU2D add_15809_17 (.A0(recv_buffer[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18601), .COUT(n18602));
    defparam add_15809_17.INIT0 = 16'hf555;
    defparam add_15809_17.INIT1 = 16'hf555;
    defparam add_15809_17.INJECT1_0 = "NO";
    defparam add_15809_17.INJECT1_1 = "NO";
    FD1P3JX speed_set_m1_i0_i19 (.D(recv_buffer[94]), .SP(clkout_c_enable_245), 
            .PD(n12617), .CK(clkout_c), .Q(speed_set_m1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i20 (.D(recv_buffer[95]), .SP(clkout_c_enable_245), 
            .CD(n12617), .CK(clkout_c), .Q(speed_set_m1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i20.GSR = "DISABLED";
    CCU2D add_15809_15 (.A0(recv_buffer[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18600), .COUT(n18601));
    defparam add_15809_15.INIT0 = 16'h0aaa;
    defparam add_15809_15.INIT1 = 16'hf555;
    defparam add_15809_15.INJECT1_0 = "NO";
    defparam add_15809_15.INJECT1_1 = "NO";
    CCU2D add_15809_13 (.A0(recv_buffer[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18599), .COUT(n18600));
    defparam add_15809_13.INIT0 = 16'hf555;
    defparam add_15809_13.INIT1 = 16'hf555;
    defparam add_15809_13.INJECT1_0 = "NO";
    defparam add_15809_13.INJECT1_1 = "NO";
    FD1P3JX speed_set_m2_i0_i1 (.D(recv_buffer[55]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i1.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i2 (.D(recv_buffer[56]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i2.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i3 (.D(recv_buffer[57]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i4 (.D(recv_buffer[58]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i4.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i5 (.D(recv_buffer[59]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i6 (.D(recv_buffer[60]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i7 (.D(recv_buffer[61]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i8 (.D(recv_buffer[62]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i9 (.D(recv_buffer[63]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i9.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i10 (.D(recv_buffer[64]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i11 (.D(recv_buffer[65]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i11.GSR = "DISABLED";
    CCU2D add_15809_11 (.A0(recv_buffer[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18598), .COUT(n18599));
    defparam add_15809_11.INIT0 = 16'h0aaa;
    defparam add_15809_11.INIT1 = 16'h0aaa;
    defparam add_15809_11.INJECT1_0 = "NO";
    defparam add_15809_11.INJECT1_1 = "NO";
    CCU2D add_15809_9 (.A0(recv_buffer[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18597), .COUT(n18598));
    defparam add_15809_9.INIT0 = 16'hf555;
    defparam add_15809_9.INIT1 = 16'h0aaa;
    defparam add_15809_9.INJECT1_0 = "NO";
    defparam add_15809_9.INJECT1_1 = "NO";
    FD1P3IX speed_set_m2_i0_i12 (.D(recv_buffer[66]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i12.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i13 (.D(recv_buffer[67]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i13.GSR = "DISABLED";
    CCU2D add_15809_7 (.A0(recv_buffer[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18596), .COUT(n18597));
    defparam add_15809_7.INIT0 = 16'hf555;
    defparam add_15809_7.INIT1 = 16'hf555;
    defparam add_15809_7.INJECT1_0 = "NO";
    defparam add_15809_7.INJECT1_1 = "NO";
    CCU2D add_15809_5 (.A0(recv_buffer[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18595), .COUT(n18596));
    defparam add_15809_5.INIT0 = 16'hf555;
    defparam add_15809_5.INIT1 = 16'h0aaa;
    defparam add_15809_5.INJECT1_0 = "NO";
    defparam add_15809_5.INJECT1_1 = "NO";
    FD1P3JX speed_set_m2_i0_i14 (.D(recv_buffer[68]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i15 (.D(recv_buffer[69]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i15.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i16 (.D(recv_buffer[70]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i16.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i17 (.D(recv_buffer[71]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i17.GSR = "DISABLED";
    CCU2D add_15803_16 (.A0(recv_buffer[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18662), .S1(n3479));
    defparam add_15803_16.INIT0 = 16'h0aaa;
    defparam add_15803_16.INIT1 = 16'h0000;
    defparam add_15803_16.INJECT1_0 = "NO";
    defparam add_15803_16.INJECT1_1 = "NO";
    FD1P3JX speed_set_m2_i0_i18 (.D(recv_buffer[72]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i18.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i19 (.D(recv_buffer[73]), .SP(clkout_c_enable_245), 
            .PD(n12597), .CK(clkout_c), .Q(speed_set_m2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i20 (.D(recv_buffer[74]), .SP(clkout_c_enable_245), 
            .CD(n12597), .CK(clkout_c), .Q(speed_set_m2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i20.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(hallsense_m2[2]), .B(n21597), .C(dir_m2), .D(hallsense_m2[1]), 
         .Z(n2915)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut.init = 16'h4008;
    FD1P3JX speed_set_m3_i0_i1 (.D(recv_buffer[34]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_129 (.A(hallsense_m2[1]), .B(n21597), .C(dir_m2), 
         .D(hallsense_m2[0]), .Z(n2951)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_129.init = 16'h4008;
    CCU2D add_15809_3 (.A0(recv_buffer[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18594), .COUT(n18595));
    defparam add_15809_3.INIT0 = 16'hf555;
    defparam add_15809_3.INIT1 = 16'hf555;
    defparam add_15809_3.INJECT1_0 = "NO";
    defparam add_15809_3.INJECT1_1 = "NO";
    FD1P3JX speed_set_m3_i0_i2 (.D(recv_buffer[35]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i2.GSR = "DISABLED";
    CCU2D add_15803_14 (.A0(recv_buffer[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18661), .COUT(n18662));
    defparam add_15803_14.INIT0 = 16'h5aaa;
    defparam add_15803_14.INIT1 = 16'h5aaa;
    defparam add_15803_14.INJECT1_0 = "NO";
    defparam add_15803_14.INJECT1_1 = "NO";
    CCU2D add_15803_12 (.A0(recv_buffer[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18660), .COUT(n18661));
    defparam add_15803_12.INIT0 = 16'h5aaa;
    defparam add_15803_12.INIT1 = 16'h5aaa;
    defparam add_15803_12.INJECT1_0 = "NO";
    defparam add_15803_12.INJECT1_1 = "NO";
    FD1P3JX speed_set_m3_i0_i3 (.D(recv_buffer[36]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i3.GSR = "DISABLED";
    CCU2D add_15803_10 (.A0(recv_buffer[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18659), .COUT(n18660));
    defparam add_15803_10.INIT0 = 16'h5555;
    defparam add_15803_10.INIT1 = 16'h5aaa;
    defparam add_15803_10.INJECT1_0 = "NO";
    defparam add_15803_10.INJECT1_1 = "NO";
    CCU2D add_15803_8 (.A0(recv_buffer[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18658), .COUT(n18659));
    defparam add_15803_8.INIT0 = 16'h5aaa;
    defparam add_15803_8.INIT1 = 16'h5aaa;
    defparam add_15803_8.INJECT1_0 = "NO";
    defparam add_15803_8.INJECT1_1 = "NO";
    FD1P3JX speed_set_m3_i0_i4 (.D(recv_buffer[37]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i4.GSR = "DISABLED";
    CCU2D add_15803_6 (.A0(recv_buffer[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18657), .COUT(n18658));
    defparam add_15803_6.INIT0 = 16'h5555;
    defparam add_15803_6.INIT1 = 16'h5555;
    defparam add_15803_6.INJECT1_0 = "NO";
    defparam add_15803_6.INJECT1_1 = "NO";
    CCU2D add_15809_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[33]), .B1(recv_buffer[34]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18594));
    defparam add_15809_1.INIT0 = 16'hF000;
    defparam add_15809_1.INIT1 = 16'ha666;
    defparam add_15809_1.INJECT1_0 = "NO";
    defparam add_15809_1.INJECT1_1 = "NO";
    FD1P3JX speed_set_m3_i0_i5 (.D(recv_buffer[38]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i6 (.D(recv_buffer[39]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i7 (.D(recv_buffer[40]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i8 (.D(recv_buffer[41]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i8.GSR = "DISABLED";
    CCU2D add_15803_4 (.A0(recv_buffer[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18656), .COUT(n18657));
    defparam add_15803_4.INIT0 = 16'h5aaa;
    defparam add_15803_4.INIT1 = 16'h5555;
    defparam add_15803_4.INJECT1_0 = "NO";
    defparam add_15803_4.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_130 (.A(hallsense_m3[2]), .B(n21592), .C(dir_m3), 
         .D(hallsense_m3[1]), .Z(n3045)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_130.init = 16'h4008;
    LUT4 i1_4_lut_adj_131 (.A(hallsense_m3[1]), .B(n21592), .C(dir_m3), 
         .D(hallsense_m3[0]), .Z(n3081)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_131.init = 16'h4008;
    LUT4 i3_4_lut (.A(SCKold), .B(n22203), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_96)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut.init = 16'h0400;
    CCU2D add_15803_2 (.A0(recv_buffer[18]), .B0(recv_buffer[17]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18656));
    defparam add_15803_2.INIT0 = 16'h7000;
    defparam add_15803_2.INIT1 = 16'h5aaa;
    defparam add_15803_2.INJECT1_0 = "NO";
    defparam add_15803_2.INJECT1_1 = "NO";
    CCU2D add_15804_21 (.A0(recv_buffer[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18655), .S1(n3455));
    defparam add_15804_21.INIT0 = 16'h5555;
    defparam add_15804_21.INIT1 = 16'h0000;
    defparam add_15804_21.INJECT1_0 = "NO";
    defparam add_15804_21.INJECT1_1 = "NO";
    CCU2D add_15804_19 (.A0(recv_buffer[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18654), .COUT(n18655));
    defparam add_15804_19.INIT0 = 16'hf555;
    defparam add_15804_19.INIT1 = 16'hf555;
    defparam add_15804_19.INJECT1_0 = "NO";
    defparam add_15804_19.INJECT1_1 = "NO";
    CCU2D add_15804_17 (.A0(recv_buffer[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18653), .COUT(n18654));
    defparam add_15804_17.INIT0 = 16'hf555;
    defparam add_15804_17.INIT1 = 16'hf555;
    defparam add_15804_17.INJECT1_0 = "NO";
    defparam add_15804_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_132 (.A(hallsense_m4[2]), .B(n21588), .C(dir_m4), 
         .D(hallsense_m4[1]), .Z(n3175)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_132.init = 16'h4008;
    LUT4 i1_4_lut_adj_133 (.A(hallsense_m4[1]), .B(n21588), .C(dir_m4), 
         .D(hallsense_m4[0]), .Z(n3211)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_133.init = 16'h4008;
    LUT4 i2_4_lut_adj_134 (.A(n3335), .B(n3311), .C(n39_adj_1894), .D(n40_adj_1895), 
         .Z(enable_m1_N_627)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_134.init = 16'h8880;
    LUT4 i18_4_lut_adj_135 (.A(recv_buffer[88]), .B(n36_adj_1896), .C(n28_adj_1897), 
         .D(recv_buffer[87]), .Z(n39_adj_1894)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i18_4_lut_adj_135.init = 16'hfffe;
    LUT4 i19_4_lut_adj_136 (.A(recv_buffer[90]), .B(n38_adj_1898), .C(n32_adj_1899), 
         .D(recv_buffer[85]), .Z(n40_adj_1895)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i19_4_lut_adj_136.init = 16'hfffe;
    LUT4 i15_4_lut_adj_137 (.A(recv_buffer[75]), .B(recv_buffer[82]), .C(recv_buffer[92]), 
         .D(recv_buffer[86]), .Z(n36_adj_1896)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i15_4_lut_adj_137.init = 16'hfffe;
    LUT4 i7_2_lut_adj_138 (.A(recv_buffer[76]), .B(recv_buffer[77]), .Z(n28_adj_1897)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i7_2_lut_adj_138.init = 16'heeee;
    LUT4 i17_4_lut_adj_139 (.A(recv_buffer[83]), .B(n34_adj_1900), .C(n24_adj_1901), 
         .D(recv_buffer[91]), .Z(n38_adj_1898)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i17_4_lut_adj_139.init = 16'hfffe;
    CCU2D add_15804_15 (.A0(recv_buffer[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18652), .COUT(n18653));
    defparam add_15804_15.INIT0 = 16'h0aaa;
    defparam add_15804_15.INIT1 = 16'hf555;
    defparam add_15804_15.INJECT1_0 = "NO";
    defparam add_15804_15.INJECT1_1 = "NO";
    LUT4 i11_3_lut_adj_140 (.A(recv_buffer[81]), .B(recv_buffer[78]), .C(recv_buffer[89]), 
         .Z(n32_adj_1899)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i11_3_lut_adj_140.init = 16'hfefe;
    LUT4 i13_4_lut_adj_141 (.A(recv_buffer[95]), .B(recv_buffer[94]), .C(recv_buffer[84]), 
         .D(recv_buffer[79]), .Z(n34_adj_1900)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i13_4_lut_adj_141.init = 16'hfffe;
    LUT4 i3_2_lut_adj_142 (.A(recv_buffer[93]), .B(recv_buffer[80]), .Z(n24_adj_1901)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(146[7:28])
    defparam i3_2_lut_adj_142.init = 16'heeee;
    CCU2D add_15804_13 (.A0(recv_buffer[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18651), .COUT(n18652));
    defparam add_15804_13.INIT0 = 16'hf555;
    defparam add_15804_13.INIT1 = 16'hf555;
    defparam add_15804_13.INJECT1_0 = "NO";
    defparam add_15804_13.INJECT1_1 = "NO";
    CCU2D add_15804_11 (.A0(recv_buffer[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18650), .COUT(n18651));
    defparam add_15804_11.INIT0 = 16'h0aaa;
    defparam add_15804_11.INIT1 = 16'h0aaa;
    defparam add_15804_11.INJECT1_0 = "NO";
    defparam add_15804_11.INJECT1_1 = "NO";
    CCU2D add_15804_9 (.A0(recv_buffer[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18649), .COUT(n18650));
    defparam add_15804_9.INIT0 = 16'hf555;
    defparam add_15804_9.INIT1 = 16'h0aaa;
    defparam add_15804_9.INJECT1_0 = "NO";
    defparam add_15804_9.INJECT1_1 = "NO";
    CCU2D add_15804_7 (.A0(recv_buffer[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18648), .COUT(n18649));
    defparam add_15804_7.INIT0 = 16'hf555;
    defparam add_15804_7.INIT1 = 16'hf555;
    defparam add_15804_7.INJECT1_0 = "NO";
    defparam add_15804_7.INJECT1_1 = "NO";
    CCU2D add_15804_5 (.A0(recv_buffer[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18647), .COUT(n18648));
    defparam add_15804_5.INIT0 = 16'hf555;
    defparam add_15804_5.INIT1 = 16'h0aaa;
    defparam add_15804_5.INJECT1_0 = "NO";
    defparam add_15804_5.INJECT1_1 = "NO";
    CCU2D add_15804_3 (.A0(recv_buffer[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18646), .COUT(n18647));
    defparam add_15804_3.INIT0 = 16'hf555;
    defparam add_15804_3.INIT1 = 16'hf555;
    defparam add_15804_3.INJECT1_0 = "NO";
    defparam add_15804_3.INJECT1_1 = "NO";
    CCU2D add_15804_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n169[0]), .B1(recv_buffer[13]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18646));
    defparam add_15804_1.INIT0 = 16'hF000;
    defparam add_15804_1.INIT1 = 16'ha666;
    defparam add_15804_1.INJECT1_0 = "NO";
    defparam add_15804_1.INJECT1_1 = "NO";
    CCU2D add_15797_21 (.A0(recv_buffer[95]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18727), .S1(n3311));
    defparam add_15797_21.INIT0 = 16'h5555;
    defparam add_15797_21.INIT1 = 16'h0000;
    defparam add_15797_21.INJECT1_0 = "NO";
    defparam add_15797_21.INJECT1_1 = "NO";
    FD1P3JX speed_set_m3_i0_i9 (.D(recv_buffer[42]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i9.GSR = "DISABLED";
    CCU2D add_15797_19 (.A0(recv_buffer[93]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[94]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18726), .COUT(n18727));
    defparam add_15797_19.INIT0 = 16'hf555;
    defparam add_15797_19.INIT1 = 16'hf555;
    defparam add_15797_19.INJECT1_0 = "NO";
    defparam add_15797_19.INJECT1_1 = "NO";
    CCU2D add_15797_17 (.A0(recv_buffer[91]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[92]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18725), .COUT(n18726));
    defparam add_15797_17.INIT0 = 16'hf555;
    defparam add_15797_17.INIT1 = 16'hf555;
    defparam add_15797_17.INJECT1_0 = "NO";
    defparam add_15797_17.INJECT1_1 = "NO";
    CCU2D add_15797_15 (.A0(recv_buffer[89]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[90]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18724), .COUT(n18725));
    defparam add_15797_15.INIT0 = 16'h0aaa;
    defparam add_15797_15.INIT1 = 16'hf555;
    defparam add_15797_15.INJECT1_0 = "NO";
    defparam add_15797_15.INJECT1_1 = "NO";
    CCU2D add_15797_13 (.A0(recv_buffer[87]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[88]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18723), .COUT(n18724));
    defparam add_15797_13.INIT0 = 16'hf555;
    defparam add_15797_13.INIT1 = 16'hf555;
    defparam add_15797_13.INJECT1_0 = "NO";
    defparam add_15797_13.INJECT1_1 = "NO";
    CCU2D add_15797_11 (.A0(recv_buffer[85]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[86]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18722), .COUT(n18723));
    defparam add_15797_11.INIT0 = 16'h0aaa;
    defparam add_15797_11.INIT1 = 16'h0aaa;
    defparam add_15797_11.INJECT1_0 = "NO";
    defparam add_15797_11.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_143 (.A(n3383), .B(n3359), .C(n39_adj_1902), .D(n40_adj_1903), 
         .Z(enable_m2_N_635)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_143.init = 16'h8880;
    LUT4 i18_4_lut_adj_144 (.A(recv_buffer[67]), .B(n36_adj_1904), .C(n28_adj_1905), 
         .D(recv_buffer[66]), .Z(n39_adj_1902)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_144.init = 16'hfffe;
    LUT4 i19_4_lut_adj_145 (.A(recv_buffer[69]), .B(n38_adj_1906), .C(n32_adj_1907), 
         .D(recv_buffer[64]), .Z(n40_adj_1903)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_145.init = 16'hfffe;
    LUT4 i15_4_lut_adj_146 (.A(recv_buffer[54]), .B(recv_buffer[61]), .C(recv_buffer[71]), 
         .D(recv_buffer[65]), .Z(n36_adj_1904)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_146.init = 16'hfffe;
    LUT4 i7_2_lut_adj_147 (.A(recv_buffer[55]), .B(recv_buffer[56]), .Z(n28_adj_1905)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_147.init = 16'heeee;
    LUT4 i17_4_lut_adj_148 (.A(recv_buffer[62]), .B(n34_adj_1908), .C(n24_adj_1909), 
         .D(recv_buffer[70]), .Z(n38_adj_1906)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_148.init = 16'hfffe;
    LUT4 i11_3_lut_adj_149 (.A(recv_buffer[60]), .B(recv_buffer[57]), .C(recv_buffer[68]), 
         .Z(n32_adj_1907)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_149.init = 16'hfefe;
    LUT4 i13_4_lut_adj_150 (.A(recv_buffer[74]), .B(recv_buffer[73]), .C(recv_buffer[63]), 
         .D(recv_buffer[58]), .Z(n34_adj_1908)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_150.init = 16'hfffe;
    LUT4 i3_2_lut_adj_151 (.A(recv_buffer[72]), .B(recv_buffer[59]), .Z(n24_adj_1909)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_151.init = 16'heeee;
    LUT4 i2_4_lut_adj_152 (.A(n3431), .B(n3407), .C(n39_adj_1910), .D(n40_adj_1911), 
         .Z(enable_m3_N_642)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_152.init = 16'h8880;
    LUT4 i18_4_lut_adj_153 (.A(recv_buffer[46]), .B(n36_adj_1912), .C(n28_adj_1913), 
         .D(recv_buffer[45]), .Z(n39_adj_1910)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_153.init = 16'hfffe;
    LUT4 i19_4_lut_adj_154 (.A(recv_buffer[48]), .B(n38_adj_1914), .C(n32_adj_1915), 
         .D(recv_buffer[43]), .Z(n40_adj_1911)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_154.init = 16'hfffe;
    LUT4 i15_4_lut_adj_155 (.A(recv_buffer[33]), .B(recv_buffer[40]), .C(recv_buffer[50]), 
         .D(recv_buffer[44]), .Z(n36_adj_1912)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_155.init = 16'hfffe;
    LUT4 i7_2_lut_adj_156 (.A(recv_buffer[34]), .B(recv_buffer[35]), .Z(n28_adj_1913)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_156.init = 16'heeee;
    LUT4 i17_4_lut_adj_157 (.A(recv_buffer[41]), .B(n34_adj_1916), .C(n24_adj_1917), 
         .D(recv_buffer[49]), .Z(n38_adj_1914)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_157.init = 16'hfffe;
    LUT4 i11_3_lut_adj_158 (.A(recv_buffer[39]), .B(recv_buffer[36]), .C(recv_buffer[47]), 
         .Z(n32_adj_1915)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_158.init = 16'hfefe;
    LUT4 i13_4_lut_adj_159 (.A(recv_buffer[53]), .B(recv_buffer[52]), .C(recv_buffer[42]), 
         .D(recv_buffer[37]), .Z(n34_adj_1916)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_159.init = 16'hfffe;
    LUT4 i3_2_lut_adj_160 (.A(recv_buffer[51]), .B(recv_buffer[38]), .Z(n24_adj_1917)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_160.init = 16'heeee;
    FD1P3IX speed_set_m3_i0_i10 (.D(recv_buffer[43]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i11 (.D(recv_buffer[44]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i12 (.D(recv_buffer[45]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i12.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i13 (.D(recv_buffer[46]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i13.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i14 (.D(recv_buffer[47]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i15 (.D(recv_buffer[48]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i15.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i16 (.D(recv_buffer[49]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i16.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i17 (.D(recv_buffer[50]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i17.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i18 (.D(recv_buffer[51]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i18.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i19 (.D(recv_buffer[52]), .SP(clkout_c_enable_245), 
            .PD(n12577), .CK(clkout_c), .Q(speed_set_m3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i20 (.D(recv_buffer[53]), .SP(clkout_c_enable_245), 
            .CD(n12577), .CK(clkout_c), .Q(speed_set_m3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i20.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i1 (.D(recv_buffer[13]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i1.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i2 (.D(recv_buffer[14]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i2.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i3 (.D(recv_buffer[15]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i4 (.D(recv_buffer[16]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i4.GSR = "DISABLED";
    CCU2D add_15797_9 (.A0(recv_buffer[83]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[84]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18721), .COUT(n18722));
    defparam add_15797_9.INIT0 = 16'hf555;
    defparam add_15797_9.INIT1 = 16'h0aaa;
    defparam add_15797_9.INJECT1_0 = "NO";
    defparam add_15797_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_161 (.A(hallsense_m1[2]), .B(n21574), .C(dir_m1), 
         .D(hallsense_m1[1]), .Z(n2785)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_161.init = 16'h4008;
    CCU2D add_15797_7 (.A0(recv_buffer[81]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[82]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18720), .COUT(n18721));
    defparam add_15797_7.INIT0 = 16'hf555;
    defparam add_15797_7.INIT1 = 16'hf555;
    defparam add_15797_7.INJECT1_0 = "NO";
    defparam add_15797_7.INJECT1_1 = "NO";
    CCU2D add_15797_5 (.A0(recv_buffer[79]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[80]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18719), .COUT(n18720));
    defparam add_15797_5.INIT0 = 16'hf555;
    defparam add_15797_5.INIT1 = 16'h0aaa;
    defparam add_15797_5.INJECT1_0 = "NO";
    defparam add_15797_5.INJECT1_1 = "NO";
    CCU2D add_15797_3 (.A0(recv_buffer[77]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[78]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18718), .COUT(n18719));
    defparam add_15797_3.INIT0 = 16'hf555;
    defparam add_15797_3.INIT1 = 16'hf555;
    defparam add_15797_3.INJECT1_0 = "NO";
    defparam add_15797_3.INJECT1_1 = "NO";
    CCU2D add_15797_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[75]), .B1(recv_buffer[76]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18718));
    defparam add_15797_1.INIT0 = 16'hF000;
    defparam add_15797_1.INIT1 = 16'ha666;
    defparam add_15797_1.INJECT1_0 = "NO";
    defparam add_15797_1.INJECT1_1 = "NO";
    FD1P3JX speed_set_m4_i0_i5 (.D(recv_buffer[17]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i5.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_162 (.A(hallsense_m1[1]), .B(n21574), .C(dir_m1), 
         .D(hallsense_m1[0]), .Z(n2821)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_162.init = 16'h4008;
    FD1P3IX speed_set_m4_i0_i6 (.D(recv_buffer[18]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i7 (.D(recv_buffer[19]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i8 (.D(recv_buffer[20]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i9 (.D(recv_buffer[21]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i9.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i10 (.D(recv_buffer[22]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i11 (.D(recv_buffer[23]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i12 (.D(recv_buffer[24]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i12.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i13 (.D(recv_buffer[25]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i13.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i14 (.D(recv_buffer[26]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i15 (.D(recv_buffer[27]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i15.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i16 (.D(recv_buffer[28]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i16.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i17 (.D(recv_buffer[29]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i17.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i18 (.D(recv_buffer[30]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i18.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i19 (.D(recv_buffer[31]), .SP(clkout_c_enable_245), 
            .PD(n12557), .CK(clkout_c), .Q(speed_set_m4[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i20 (.D(recv_buffer[32]), .SP(clkout_c_enable_245), 
            .CD(n12557), .CK(clkout_c), .Q(speed_set_m4[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=293, LSE_RLINE=293 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i20.GSR = "DISABLED";
    PFUMX i18136 (.BLUT(n21481), .ALUT(n21480), .C0(n22203), .Z(MISO_N_670));
    LUT4 SCKold_I_0_2_lut_rep_371 (.A(SCKold), .B(SCKlatched), .Z(n21580)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(193[8:45])
    defparam SCKold_I_0_2_lut_rep_371.init = 16'h2222;
    LUT4 CSlatched_I_0_1_lut_rep_372 (.A(CSlatched), .Z(n21581)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam CSlatched_I_0_1_lut_rep_372.init = 16'h5555;
    LUT4 mux_9_i24_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[23]), .C(\speed_m4[11] ), 
         .D(n22202), .Z(MISOb_N_666[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i160_2_lut_rep_347_3_lut_3_lut (.A(n22201), .B(SCKlatched), .C(SCKold), 
         .Z(n21556)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam i160_2_lut_rep_347_3_lut_3_lut.init = 16'h1010;
    LUT4 CSold_I_0_2_lut_rep_346_2_lut (.A(n22201), .B(n22202), .Z(n21555)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam CSold_I_0_2_lut_rep_346_2_lut.init = 16'h4444;
    LUT4 mux_9_i26_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[25]), .C(\speed_m4[13] ), 
         .D(n22202), .Z(MISOb_N_666[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i27_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[26]), .C(\speed_m4[14] ), 
         .D(n22202), .Z(MISOb_N_666[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i22_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[21]), .C(\speed_m4[9] ), 
         .D(n22202), .Z(MISOb_N_666[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i28_3_lut_4_lut_4_lut (.A(n22201), .B(send_buffer[27]), .C(\speed_m4[15] ), 
         .D(n22202), .Z(MISOb_N_666[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    
endmodule
//
// Verilog Description of module HALL_U4
//

module HALL_U4 (clk_1mhz, \speed_m2[0] , hallsense_m2, clkout_c_enable_176, 
            clkout_c_enable_164, H_C_m2_c, H_B_m2_c, H_A_m2_c, \speed_m2[1] , 
            \speed_m2[2] , \speed_m2[3] , \speed_m2[4] , \speed_m2[5] , 
            \speed_m2[6] , \speed_m2[7] , \speed_m2[8] , \speed_m2[9] , 
            \speed_m2[10] , \speed_m2[11] , \speed_m2[12] , \speed_m2[13] , 
            \speed_m2[14] , \speed_m2[15] , \speed_m2[16] , \speed_m2[17] , 
            \speed_m2[18] , \speed_m2[19] , GND_net, n22198);
    input clk_1mhz;
    output \speed_m2[0] ;
    output [2:0]hallsense_m2;
    input clkout_c_enable_176;
    input clkout_c_enable_164;
    input H_C_m2_c;
    input H_B_m2_c;
    input H_A_m2_c;
    output \speed_m2[1] ;
    output \speed_m2[2] ;
    output \speed_m2[3] ;
    output \speed_m2[4] ;
    output \speed_m2[5] ;
    output \speed_m2[6] ;
    output \speed_m2[7] ;
    output \speed_m2[8] ;
    output \speed_m2[9] ;
    output \speed_m2[10] ;
    output \speed_m2[11] ;
    output \speed_m2[12] ;
    output \speed_m2[13] ;
    output \speed_m2[14] ;
    output \speed_m2[15] ;
    output \speed_m2[16] ;
    output \speed_m2[17] ;
    output \speed_m2[18] ;
    output \speed_m2[19] ;
    input GND_net;
    input n22198;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(62[10:22])
    
    wire stable_counting, n21514, n21534;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_lat, hall3_old, hall1_old, hall1_lat, hall2_lat;
    wire [19:0]speedt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_85, n4333;
    wire [19:0]n7;
    
    wire hall2_old, n21760, n21761, stable_counting_N_1746, n21128, 
        n19642, n19845, n21513, n21127;
    wire [6:0]stable_counting_N_1759;
    
    wire n21533, n21532, stable_counting_N_1758, n21539, n21582, n21558;
    wire [6:0]n83;
    wire [19:0]count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(60[10:15])
    
    wire n4, n19963, n18466, n18465, n18464, n18463, n18462, n18461, 
        n18460, n18459, n18458, n18457, n19666, n10_adj_1881, n19906, 
        n12_adj_1882, n15_adj_1883, n14_adj_1884, n101, n19959, n19910, 
        n16_adj_1885, n95;
    
    FD1P3IX stable_count__i0 (.D(n21534), .SP(stable_counting), .CD(n21514), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall3_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall1_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m2_c), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall3_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m2_c), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall2_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3IX speedt__i0 (.D(n7[0]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall2_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m2_c), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall1_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    LUT4 stable_count_2__bdd_4_lut_18277 (.A(stable_count[2]), .B(stable_count[1]), 
         .C(stable_count[3]), .D(stable_count[4]), .Z(n21760)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam stable_count_2__bdd_4_lut_18277.init = 16'h7ffe;
    LUT4 i17012_4_lut_4_lut (.A(n21761), .B(stable_counting_N_1746), .C(n21128), 
         .D(n19642), .Z(n19845)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17012_4_lut_4_lut.init = 16'hfffe;
    LUT4 n12547_bdd_4_lut (.A(stable_counting_N_1746), .B(stable_count[6]), 
         .C(stable_count[5]), .D(n21513), .Z(n21127)) /* synthesis lut_function=(!(A+(B (C (D))+!B !(C+(D))))) */ ;
    defparam n12547_bdd_4_lut.init = 16'h1554;
    LUT4 i13813_2_lut_4_lut (.A(stable_count[6]), .B(stable_count[5]), .C(n21513), 
         .D(stable_counting_N_1746), .Z(stable_counting_N_1759[6])) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (((D)+!C)+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13813_2_lut_4_lut.init = 16'h006a;
    FD1P3IX stable_count__i1 (.D(stable_counting_N_1759[1]), .SP(stable_counting), 
            .CD(n21514), .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(stable_counting_N_1759[2]), .SP(stable_counting), 
            .CD(n21514), .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n21533), .SP(stable_counting), .CD(n21514), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(stable_counting_N_1759[4]), .SP(stable_counting), 
            .CD(n21514), .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(stable_counting_N_1759[5]), .SP(stable_counting), 
            .CD(n21514), .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i6 (.D(stable_counting_N_1759[6]), .SP(stable_counting), 
            .CD(n21514), .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    LUT4 i13812_2_lut_3_lut_4_lut (.A(stable_count[4]), .B(n21532), .C(stable_counting_N_1746), 
         .D(stable_count[5]), .Z(stable_counting_N_1759[5])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13812_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i2194_2_lut_rep_305 (.A(stable_counting), .B(stable_counting_N_1758), 
         .Z(n21514)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i2194_2_lut_rep_305.init = 16'h8888;
    LUT4 i17872_2_lut_rep_289_2_lut_3_lut (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21539), .Z(clk_1mhz_enable_85)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i17872_2_lut_rep_289_2_lut_3_lut.init = 16'h8f8f;
    LUT4 n780_bdd_2_lut_18019_3_lut_3_lut_4_lut (.A(stable_counting), .B(stable_counting_N_1758), 
         .C(n21127), .D(n21539), .Z(n21128)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C+(D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam n780_bdd_2_lut_18019_3_lut_3_lut_4_lut.init = 16'hf7f0;
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i2363_2_lut_rep_373 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21582)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2363_2_lut_rep_373.init = 16'h8888;
    LUT4 i2370_2_lut_rep_349_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21558)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2370_2_lut_rep_349_3_lut.init = 16'h8080;
    LUT4 i2368_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n83[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2368_2_lut_3_lut.init = 16'h7878;
    LUT4 i2377_2_lut_rep_323_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21532)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2377_2_lut_rep_323_3_lut_4_lut.init = 16'h8000;
    FD1S3IX count__i1 (.D(n7[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n7[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n7[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n7[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n7[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n7[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n7[7]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n7[8]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n7[9]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n7[10]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n7[11]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n7[12]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n7[13]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n7[14]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n7[15]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n7[16]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n7[17]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n7[18]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n7[19]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    LUT4 mux_28_i2_4_lut (.A(n7[1]), .B(speedt[1]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hac0a;
    LUT4 mux_28_i3_4_lut (.A(n7[2]), .B(speedt[2]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hac0a;
    LUT4 mux_28_i4_4_lut (.A(n7[3]), .B(speedt[3]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hac0a;
    LUT4 mux_28_i5_4_lut (.A(n7[4]), .B(speedt[4]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hac0a;
    LUT4 mux_28_i6_4_lut (.A(n7[5]), .B(speedt[5]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hac0a;
    LUT4 mux_28_i7_4_lut (.A(n7[6]), .B(speedt[6]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hac0a;
    LUT4 mux_28_i8_4_lut (.A(n7[7]), .B(speedt[7]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hac0a;
    LUT4 mux_28_i9_4_lut (.A(n7[8]), .B(speedt[8]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hac0a;
    LUT4 mux_28_i10_4_lut (.A(n7[9]), .B(speedt[9]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hac0a;
    LUT4 mux_28_i11_4_lut (.A(n7[10]), .B(speedt[10]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hac0a;
    FD1P3IX speedt__i1 (.D(n7[1]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    LUT4 mux_28_i12_4_lut (.A(n7[11]), .B(speedt[11]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hac0a;
    LUT4 mux_28_i13_4_lut (.A(n7[12]), .B(speedt[12]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hac0a;
    LUT4 mux_28_i14_4_lut (.A(n7[13]), .B(speedt[13]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hac0a;
    LUT4 mux_28_i15_4_lut (.A(n7[14]), .B(speedt[14]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hac0a;
    LUT4 mux_28_i16_4_lut (.A(n7[15]), .B(speedt[15]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hac0a;
    LUT4 i2_3_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(92[7:87])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 mux_28_i17_4_lut (.A(n7[16]), .B(speedt[16]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hac0a;
    LUT4 i17129_3_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(stable_counting_N_1758), .Z(n19963)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i17129_3_lut.init = 16'hc8c8;
    LUT4 mux_28_i18_4_lut (.A(n7[17]), .B(speedt[17]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hac0a;
    LUT4 mux_28_i19_4_lut (.A(n7[18]), .B(speedt[18]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hac0a;
    LUT4 mux_28_i20_4_lut (.A(n7[19]), .B(speedt[19]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hac0a;
    FD1P3IX speedt__i2 (.D(n7[2]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n7[3]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n7[4]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n7[5]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n7[6]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n7[7]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n7[8]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n7[9]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n7[10]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n7[11]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n7[12]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n7[13]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n7[14]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n7[15]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n7[16]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n7[17]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n7[18]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n7[19]), .SP(clk_1mhz_enable_85), .CD(n4333), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18466), 
          .S0(n7[19]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18465), .COUT(n18466), .S0(n7[17]), .S1(n7[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18464), .COUT(n18465), .S0(n7[15]), .S1(n7[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18463), .COUT(n18464), .S0(n7[13]), .S1(n7[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18462), .COUT(n18463), .S0(n7[11]), .S1(n7[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18461), .COUT(n18462), .S0(n7[9]), .S1(n7[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18460), 
          .COUT(n18461), .S0(n7[7]), .S1(n7[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    LUT4 n780_bdd_2_lut_18156 (.A(n21760), .B(stable_count[0]), .Z(n21761)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n780_bdd_2_lut_18156.init = 16'hbbbb;
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18459), 
          .COUT(n18460), .S0(n7[5]), .S1(n7[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18458), 
          .COUT(n18459), .S0(n7[3]), .S1(n7[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18457), 
          .COUT(n18458), .S0(n7[1]), .S1(n7[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18457), 
          .S1(n7[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i13811_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21558), .C(stable_counting_N_1746), 
         .D(stable_count[4]), .Z(stable_counting_N_1759[4])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13811_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i1_4_lut_rep_330 (.A(n19666), .B(n10_adj_1881), .C(n19642), .D(n19906), 
         .Z(n21539)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_4_lut_rep_330.init = 16'hf7ff;
    LUT4 mux_28_i1_4_lut (.A(n7[0]), .B(speedt[0]), .C(stable_counting_N_1758), 
         .D(n21539), .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hac0a;
    LUT4 i17072_2_lut (.A(count[1]), .B(count[5]), .Z(n19906)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17072_2_lut.init = 16'h8888;
    LUT4 i6_4_lut (.A(count[17]), .B(n12_adj_1882), .C(count[16]), .D(count[19]), 
         .Z(n19666)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[9]), .B(count[4]), .C(count[18]), .D(count[14]), 
         .Z(n12_adj_1882)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(count[3]), .B(count[2]), .Z(n10_adj_1881)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i8_4_lut (.A(n15_adj_1883), .B(count[12]), .C(n14_adj_1884), 
         .D(count[11]), .Z(n19642)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut_adj_125 (.A(count[0]), .B(count[10]), .C(count[7]), 
         .D(count[8]), .Z(n15_adj_1883)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_125.init = 16'hfffe;
    LUT4 i5_3_lut (.A(count[13]), .B(count[15]), .C(count[6]), .Z(n14_adj_1884)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut (.A(stable_count[0]), .B(n101), .C(n19959), .D(n19910), 
         .Z(stable_counting_N_1758)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[7:23])
    defparam i1_4_lut.init = 16'h0008;
    LUT4 i8_4_lut_adj_126 (.A(n19845), .B(n16_adj_1885), .C(count[5]), 
         .D(stable_counting), .Z(n4333)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i8_4_lut_adj_126.init = 16'h4000;
    LUT4 i7_4_lut (.A(n83[1]), .B(n19666), .C(count[1]), .D(n10_adj_1881), 
         .Z(n16_adj_1885)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i1_3_lut (.A(n95), .B(hall2_lat), .C(hall2_old), .Z(n101)) /* synthesis lut_function=(A (B (C)+!B !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[7:23])
    defparam i1_3_lut.init = 16'h8282;
    LUT4 i17125_4_lut (.A(stable_count[3]), .B(stable_count[5]), .C(stable_count[4]), 
         .D(stable_count[6]), .Z(n19959)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17125_4_lut.init = 16'hfffe;
    LUT4 i17962_2_lut_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), 
         .D(n83[1]), .Z(stable_counting_N_1759[1])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i17962_2_lut_2_lut_4_lut.init = 16'h2100;
    LUT4 i17854_2_lut_rep_325_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), 
         .D(stable_count[0]), .Z(n21534)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C+(D))))) */ ;
    defparam i17854_2_lut_rep_325_4_lut.init = 16'h0021;
    LUT4 i13809_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .D(n83[2]), 
         .Z(stable_counting_N_1759[2])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i13809_2_lut_4_lut.init = 16'h2100;
    LUT4 i17076_2_lut (.A(stable_count[2]), .B(stable_count[1]), .Z(n19910)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17076_2_lut.init = 16'heeee;
    LUT4 i2361_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n83[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2361_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_127 (.A(hall3_lat), .B(hall1_lat), .C(hall3_old), 
         .D(hall1_old), .Z(n95)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[7:23])
    defparam i1_4_lut_adj_127.init = 16'h8421;
    LUT4 i2384_2_lut_rep_304_3_lut_4_lut (.A(stable_count[2]), .B(n21582), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21513)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2384_2_lut_rep_304_3_lut_4_lut.init = 16'h8000;
    LUT4 i13810_3_lut_rep_324_4_lut (.A(stable_count[2]), .B(n21582), .C(stable_counting_N_1746), 
         .D(stable_count[3]), .Z(n21533)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13810_3_lut_rep_324_4_lut.init = 16'h0708;
    LUT4 i1_4_lut_adj_128 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_128.init = 16'h7bde;
    FD1S3IX count__i0 (.D(n7[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_85), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22198), .SP(stable_counting_N_1746), 
            .CD(n19963), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=312, LSE_RLINE=312 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module HALL_U3
//

module HALL_U3 (clk_1mhz, \speed_m3[0] , hallsense_m3, clkout_c_enable_176, 
            H_A_m3_c, H_B_m3_c, H_C_m3_c, clkout_c_enable_164, \speed_m3[1] , 
            \speed_m3[2] , \speed_m3[3] , \speed_m3[4] , \speed_m3[5] , 
            \speed_m3[6] , \speed_m3[7] , \speed_m3[8] , \speed_m3[9] , 
            \speed_m3[10] , \speed_m3[11] , \speed_m3[12] , \speed_m3[13] , 
            \speed_m3[14] , \speed_m3[15] , \speed_m3[16] , \speed_m3[17] , 
            \speed_m3[18] , \speed_m3[19] , GND_net, n22198);
    input clk_1mhz;
    output \speed_m3[0] ;
    output [2:0]hallsense_m3;
    input clkout_c_enable_176;
    input H_A_m3_c;
    input H_B_m3_c;
    input H_C_m3_c;
    input clkout_c_enable_164;
    output \speed_m3[1] ;
    output \speed_m3[2] ;
    output \speed_m3[3] ;
    output \speed_m3[4] ;
    output \speed_m3[5] ;
    output \speed_m3[6] ;
    output \speed_m3[7] ;
    output \speed_m3[8] ;
    output \speed_m3[9] ;
    output \speed_m3[10] ;
    output \speed_m3[11] ;
    output \speed_m3[12] ;
    output \speed_m3[13] ;
    output \speed_m3[14] ;
    output \speed_m3[15] ;
    output \speed_m3[16] ;
    output \speed_m3[17] ;
    output \speed_m3[18] ;
    output \speed_m3[19] ;
    input GND_net;
    input n22198;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(62[10:22])
    
    wire stable_counting, n21493, n21538;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_lat, hall1_lat, hall2_lat, hall3_old, hall1_old, hall2_old;
    wire [19:0]speedt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_104, n4331;
    wire [19:0]n7;
    
    wire stable_counting_N_1758, n21502, n21501;
    wire [19:0]count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(60[10:15])
    
    wire stable_counting_N_1746, n19813, n21515, n21516;
    wire [6:0]stable_counting_N_1759;
    
    wire n19999, n22, n17, n14, n18951, n19891, n22_adj_1872, 
        n21536, n21496, n21531, n19961, n13_adj_1876, n21594, n21559, 
        n18476, n21537, n18475, n21560, n16242, n18474, n18473, 
        n18472, n18471, n18470, n18469, n18468, n18467, n4, n19991, 
        n21517, n19821, n18_adj_1877, n15_adj_1878, n11_adj_1879, 
        n20_adj_1880, n19987, n19947;
    
    FD1P3IX stable_count__i0 (.D(n21538), .SP(stable_counting), .CD(n21493), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m3_c), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall1_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m3_c), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall2_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m3_c), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall3_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall3_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall1_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall2_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3IX speedt__i0 (.D(n7[0]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    LUT4 i2198_2_lut_rep_284 (.A(stable_counting), .B(stable_counting_N_1758), 
         .Z(n21493)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i2198_2_lut_rep_284.init = 16'h8888;
    LUT4 i16981_3_lut_4_lut (.A(n21502), .B(n21501), .C(count[8]), .D(stable_counting_N_1746), 
         .Z(n19813)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;
    defparam i16981_3_lut_4_lut.init = 16'hf0fe;
    LUT4 i17869_2_lut_3_lut_3_lut (.A(n21515), .B(stable_counting_N_1758), 
         .C(stable_counting), .Z(clk_1mhz_enable_104)) /* synthesis lut_function=((B (C))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i17869_2_lut_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i13846_2_lut_4_lut (.A(stable_count[6]), .B(stable_count[5]), .C(n21516), 
         .D(stable_counting_N_1746), .Z(stable_counting_N_1759[6])) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (((D)+!C)+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13846_2_lut_4_lut.init = 16'h006a;
    LUT4 i11_4_lut_4_lut (.A(n21538), .B(n19999), .C(n22), .D(n17), 
         .Z(n4331)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i11_4_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_rep_306 (.A(n14), .B(n18951), .C(n19891), .D(n22_adj_1872), 
         .Z(n21515)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_4_lut_rep_306.init = 16'hdfff;
    LUT4 i13845_2_lut_3_lut_4_lut (.A(stable_count[4]), .B(n21536), .C(stable_counting_N_1746), 
         .D(stable_count[5]), .Z(stable_counting_N_1759[5])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13845_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i2446_3_lut_rep_292_4_lut (.A(stable_count[4]), .B(n21536), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n21501)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2446_3_lut_rep_292_4_lut.init = 16'h7f80;
    LUT4 i14095_2_lut_rep_287_4_lut_3_lut_4_lut (.A(stable_count[4]), .B(n21536), 
         .C(stable_count[6]), .D(stable_count[5]), .Z(n21496)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i14095_2_lut_rep_287_4_lut_3_lut_4_lut.init = 16'h7ff8;
    FD1P3IX stable_count__i1 (.D(n21531), .SP(stable_counting), .CD(n21493), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(stable_counting_N_1759[2]), .SP(stable_counting), 
            .CD(n21493), .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(stable_counting_N_1759[3]), .SP(stable_counting), 
            .CD(n21493), .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(stable_counting_N_1759[4]), .SP(stable_counting), 
            .CD(n21493), .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(stable_counting_N_1759[5]), .SP(stable_counting), 
            .CD(n21493), .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i6 (.D(stable_counting_N_1759[6]), .SP(stable_counting), 
            .CD(n21493), .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n7[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n7[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n7[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n7[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n7[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n7[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n7[7]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n7[8]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n7[9]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n7[10]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n7[11]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n7[12]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n7[13]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n7[14]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n7[15]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n7[16]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n7[17]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n7[18]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n7[19]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i17127_3_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(stable_counting_N_1758), .Z(n19961)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i17127_3_lut.init = 16'hc8c8;
    LUT4 i17057_3_lut_4_lut (.A(count[17]), .B(count[16]), .C(count[9]), 
         .D(count[14]), .Z(n19891)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i17057_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_28_i2_4_lut (.A(n7[1]), .B(speedt[1]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hac0a;
    LUT4 mux_28_i3_4_lut (.A(n7[2]), .B(speedt[2]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hac0a;
    LUT4 i1_2_lut_3_lut (.A(count[17]), .B(count[16]), .C(n14), .Z(n13_adj_1876)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i2413_2_lut_rep_385 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21594)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2413_2_lut_rep_385.init = 16'h8888;
    LUT4 i2420_2_lut_rep_350_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21559)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2420_2_lut_rep_350_3_lut.init = 16'h8080;
    LUT4 mux_28_i4_4_lut (.A(n7[3]), .B(speedt[3]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hac0a;
    LUT4 mux_28_i5_4_lut (.A(n7[4]), .B(speedt[4]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hac0a;
    LUT4 mux_28_i6_4_lut (.A(n7[5]), .B(speedt[5]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hac0a;
    LUT4 mux_28_i7_4_lut (.A(n7[6]), .B(speedt[6]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hac0a;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18476), 
          .S0(n7[19]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    LUT4 i2427_2_lut_rep_327_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21536)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2427_2_lut_rep_327_3_lut_4_lut.init = 16'h8000;
    LUT4 i2425_2_lut_rep_328_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21537)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2425_2_lut_rep_328_3_lut_4_lut.init = 16'h78f0;
    LUT4 i13842_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_counting_N_1746), .D(stable_count[2]), .Z(stable_counting_N_1759[2])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13842_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 mux_28_i8_4_lut (.A(n7[7]), .B(speedt[7]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hac0a;
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18475), .COUT(n18476), .S0(n7[17]), .S1(n7[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    LUT4 mux_28_i9_4_lut (.A(n7[8]), .B(speedt[8]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hac0a;
    FD1P3IX speedt__i1 (.D(n7[1]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    LUT4 i2418_2_lut_rep_351_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21560)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2418_2_lut_rep_351_3_lut.init = 16'h7878;
    LUT4 mux_28_i10_4_lut (.A(n7[9]), .B(speedt[9]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hac0a;
    LUT4 mux_28_i11_4_lut (.A(n7[10]), .B(speedt[10]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hac0a;
    LUT4 mux_28_i12_4_lut (.A(n7[11]), .B(speedt[11]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hac0a;
    LUT4 mux_28_i13_4_lut (.A(n7[12]), .B(speedt[12]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hac0a;
    LUT4 mux_28_i14_4_lut (.A(n7[13]), .B(speedt[13]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hac0a;
    LUT4 mux_28_i15_4_lut (.A(n7[14]), .B(speedt[14]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hac0a;
    FD1P3IX speedt__i2 (.D(n7[2]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n7[3]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n7[4]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n7[5]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n7[6]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n7[7]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n7[8]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n7[9]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n7[10]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n7[11]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n7[12]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n7[13]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n7[14]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n7[15]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n7[16]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n7[17]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n7[18]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n7[19]), .SP(clk_1mhz_enable_104), .CD(n4331), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    LUT4 mux_28_i16_4_lut (.A(n7[15]), .B(speedt[15]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hac0a;
    LUT4 i1_2_lut_3_lut_4_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n16242)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i1_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h7ff8;
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18474), .COUT(n18475), .S0(n7[15]), .S1(n7[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18473), .COUT(n18474), .S0(n7[13]), .S1(n7[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    LUT4 mux_28_i17_4_lut (.A(n7[16]), .B(speedt[16]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hac0a;
    LUT4 mux_28_i18_4_lut (.A(n7[17]), .B(speedt[17]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hac0a;
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18472), .COUT(n18473), .S0(n7[11]), .S1(n7[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18471), .COUT(n18472), .S0(n7[9]), .S1(n7[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    LUT4 mux_28_i19_4_lut (.A(n7[18]), .B(speedt[18]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hac0a;
    LUT4 mux_28_i20_4_lut (.A(n7[19]), .B(speedt[19]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hac0a;
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18470), 
          .COUT(n18471), .S0(n7[7]), .S1(n7[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18469), 
          .COUT(n18470), .S0(n7[5]), .S1(n7[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18468), 
          .COUT(n18469), .S0(n7[3]), .S1(n7[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18467), 
          .COUT(n18468), .S0(n7[1]), .S1(n7[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18467), 
          .S1(n7[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i13841_3_lut_rep_322 (.A(stable_count[1]), .B(stable_counting_N_1746), 
         .C(stable_count[0]), .Z(n21531)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(98[4] 103[11])
    defparam i13841_3_lut_rep_322.init = 16'h1212;
    LUT4 i5_2_lut_4_lut (.A(stable_count[1]), .B(stable_counting_N_1746), 
         .C(stable_count[0]), .D(count[19]), .Z(n17)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(98[4] 103[11])
    defparam i5_2_lut_4_lut.init = 16'h1200;
    LUT4 i2439_2_lut_rep_293_3_lut_4_lut (.A(stable_count[3]), .B(n21559), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21502)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2439_2_lut_rep_293_3_lut_4_lut.init = 16'h78f0;
    LUT4 i13844_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21559), .C(stable_counting_N_1746), 
         .D(stable_count[4]), .Z(stable_counting_N_1759[4])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13844_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i1_4_lut (.A(hall2_old), .B(hall1_old), .C(hall2_lat), .D(hall1_lat), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i3_4_lut (.A(stable_count[0]), .B(stable_counting_N_1746), .C(stable_count[1]), 
         .D(n19991), .Z(stable_counting_N_1758)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[7:23])
    defparam i3_4_lut.init = 16'h0002;
    LUT4 i17157_4_lut (.A(n21496), .B(n21560), .C(n21537), .D(n21517), 
         .Z(n19991)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17157_4_lut.init = 16'hfffe;
    LUT4 mux_28_i1_4_lut (.A(n7[0]), .B(speedt[0]), .C(stable_counting_N_1758), 
         .D(n21515), .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hac0a;
    LUT4 i9_4_lut (.A(n19821), .B(n18_adj_1877), .C(count[8]), .D(count[0]), 
         .Z(n18951)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i42_2_lut (.A(count[5]), .B(count[2]), .Z(n22_adj_1872)) /* synthesis lut_function=(A (B)) */ ;
    defparam i42_2_lut.init = 16'h8888;
    LUT4 i8_4_lut (.A(n15_adj_1878), .B(n11_adj_1879), .C(count[19]), 
         .D(count[12]), .Z(n18_adj_1877)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i8_4_lut.init = 16'hffef;
    LUT4 i5_2_lut (.A(count[15]), .B(count[13]), .Z(n15_adj_1878)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(count[11]), .B(count[6]), .Z(n11_adj_1879)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i16989_2_lut (.A(count[10]), .B(count[7]), .Z(n19821)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16989_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_123 (.A(count[4]), .B(count[1]), .C(count[18]), 
         .D(count[3]), .Z(n14)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_123.init = 16'h8000;
    LUT4 i2434_2_lut_rep_307_3_lut_4_lut (.A(stable_count[2]), .B(n21594), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21516)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2434_2_lut_rep_307_3_lut_4_lut.init = 16'h8000;
    LUT4 i2432_2_lut_rep_308_3_lut_4_lut (.A(stable_count[2]), .B(n21594), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21517)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2432_2_lut_rep_308_3_lut_4_lut.init = 16'h78f0;
    LUT4 i13843_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21594), .C(stable_counting_N_1746), 
         .D(stable_count[3]), .Z(stable_counting_N_1759[3])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13843_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i10_4_lut (.A(n13_adj_1876), .B(n20_adj_1880), .C(count[5]), 
         .D(clk_1mhz_enable_104), .Z(n22)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i10_4_lut.init = 16'h8000;
    LUT4 i17165_4_lut (.A(count[13]), .B(n19987), .C(n19813), .D(count[12]), 
         .Z(n19999)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17165_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_352 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_352.init = 16'hdede;
    LUT4 i8_4_lut_adj_124 (.A(count[14]), .B(stable_counting), .C(count[2]), 
         .D(count[9]), .Z(n20_adj_1880)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut_adj_124.init = 16'h8000;
    LUT4 i17864_2_lut_rep_329_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), 
         .D(stable_count[0]), .Z(n21538)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C+(D))))) */ ;
    defparam i17864_2_lut_rep_329_4_lut.init = 16'h0021;
    LUT4 i17153_4_lut (.A(stable_counting_N_1759[4]), .B(n19947), .C(n19821), 
         .D(count[0]), .Z(n19987)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17153_4_lut.init = 16'hfffe;
    LUT4 i17113_4_lut (.A(n11_adj_1879), .B(stable_counting_N_1746), .C(count[15]), 
         .D(n16242), .Z(n19947)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i17113_4_lut.init = 16'hfbfa;
    FD1S3IX count__i0 (.D(n7[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_104), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22198), .SP(stable_counting_N_1746), 
            .CD(n19961), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module HALL_U5
//

module HALL_U5 (clk_1mhz, \speed_m1[0] , hallsense_m1, clkout_c_enable_164, 
            clkout_c_enable_176, H_A_m1_c, H_B_m1_c, H_C_m1_c, \speed_m1[1] , 
            \speed_m1[2] , \speed_m1[3] , \speed_m1[4] , \speed_m1[5] , 
            \speed_m1[6] , \speed_m1[7] , \speed_m1[8] , \speed_m1[9] , 
            \speed_m1[10] , \speed_m1[11] , \speed_m1[12] , \speed_m1[13] , 
            \speed_m1[14] , \speed_m1[15] , \speed_m1[16] , \speed_m1[17] , 
            \speed_m1[18] , \speed_m1[19] , GND_net, n22198);
    input clk_1mhz;
    output \speed_m1[0] ;
    output [2:0]hallsense_m1;
    input clkout_c_enable_164;
    input clkout_c_enable_176;
    input H_A_m1_c;
    input H_B_m1_c;
    input H_C_m1_c;
    output \speed_m1[1] ;
    output \speed_m1[2] ;
    output \speed_m1[3] ;
    output \speed_m1[4] ;
    output \speed_m1[5] ;
    output \speed_m1[6] ;
    output \speed_m1[7] ;
    output \speed_m1[8] ;
    output \speed_m1[9] ;
    output \speed_m1[10] ;
    output \speed_m1[11] ;
    output \speed_m1[12] ;
    output \speed_m1[13] ;
    output \speed_m1[14] ;
    output \speed_m1[15] ;
    output \speed_m1[16] ;
    output \speed_m1[17] ;
    output \speed_m1[18] ;
    output \speed_m1[19] ;
    input GND_net;
    input n22198;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(62[10:22])
    
    wire stable_counting, n21494, n21547;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_lat;
    wire [19:0]speedt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_66, n4298;
    wire [19:0]n7;
    
    wire hall1_old, hall1_lat, hall2_old, hall2_lat, hall3_old, n4, 
        stable_counting_N_1758, stable_counting_N_1746, n19983, n21497, 
        n21567, n21546, n21523, n21506, n21505;
    wire [19:0]count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(60[10:15])
    
    wire n19831, n21511;
    wire [6:0]stable_counting_N_1759;
    
    wire n21521, n21535, n14, n18946, n19879, n22, n20001, n22_adj_1862, 
        n17, n21545, n19965, n21606, n21566, n16318, n18456, n18455, 
        n18454, n18453, n18452, n18451, n13_adj_1866, n20_adj_1867, 
        n19989, n19953, n13_adj_1868, n11_adj_1869, n18450, n18449, 
        n18448, n18447, n18_adj_1870, n15_adj_1871;
    
    FD1P3IX stable_count__i0 (.D(n21547), .SP(stable_counting), .CD(n21494), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3IX speedt__i0 (.D(n7[0]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall1_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall2_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall3_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m1_c), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall1_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m1_c), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall2_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m1_c), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall3_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    LUT4 i17851_2_lut_rep_338_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), 
         .D(stable_count[0]), .Z(n21547)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C+(D))))) */ ;
    defparam i17851_2_lut_rep_338_4_lut.init = 16'h0021;
    LUT4 i2190_2_lut_rep_285 (.A(stable_counting), .B(stable_counting_N_1758), 
         .Z(n21494)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i2190_2_lut_rep_285.init = 16'h8888;
    LUT4 i3_4_lut (.A(stable_count[0]), .B(stable_counting_N_1746), .C(stable_count[1]), 
         .D(n19983), .Z(stable_counting_N_1758)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[7:23])
    defparam i3_4_lut.init = 16'h0002;
    LUT4 i17149_4_lut (.A(n21497), .B(n21567), .C(n21546), .D(n21523), 
         .Z(n19983)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17149_4_lut.init = 16'hfffe;
    LUT4 i16998_3_lut_4_lut (.A(n21506), .B(n21505), .C(count[8]), .D(stable_counting_N_1746), 
         .Z(n19831)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;
    defparam i16998_3_lut_4_lut.init = 16'hf0fe;
    LUT4 i17882_2_lut_3_lut_3_lut (.A(n21511), .B(stable_counting_N_1758), 
         .C(stable_counting), .Z(clk_1mhz_enable_66)) /* synthesis lut_function=((B (C))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i17882_2_lut_3_lut_3_lut.init = 16'hd5d5;
    FD1P3IX stable_count__i6 (.D(stable_counting_N_1759[6]), .SP(stable_counting), 
            .CD(n21494), .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    LUT4 i13780_2_lut_4_lut (.A(stable_count[6]), .B(stable_count[5]), .C(n21521), 
         .D(stable_counting_N_1746), .Z(stable_counting_N_1759[6])) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (((D)+!C)+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13780_2_lut_4_lut.init = 16'h006a;
    FD1P3IX stable_count__i5 (.D(stable_counting_N_1759[5]), .SP(stable_counting), 
            .CD(n21494), .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(stable_counting_N_1759[4]), .SP(stable_counting), 
            .CD(n21494), .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(stable_counting_N_1759[3]), .SP(stable_counting), 
            .CD(n21494), .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(stable_counting_N_1759[2]), .SP(stable_counting), 
            .CD(n21494), .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n21535), .SP(stable_counting), .CD(n21494), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i1_4_lut_rep_302 (.A(n14), .B(n18946), .C(n19879), .D(n22), 
         .Z(n21511)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_4_lut_rep_302.init = 16'hdfff;
    LUT4 mux_28_i2_4_lut (.A(n7[1]), .B(speedt[1]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hac0a;
    LUT4 mux_28_i3_4_lut (.A(n7[2]), .B(speedt[2]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hac0a;
    LUT4 i11_4_lut_4_lut (.A(n21547), .B(n20001), .C(n22_adj_1862), .D(n17), 
         .Z(n4298)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i11_4_lut_4_lut.init = 16'h1000;
    LUT4 mux_28_i4_4_lut (.A(n7[3]), .B(speedt[3]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hac0a;
    LUT4 mux_28_i5_4_lut (.A(n7[4]), .B(speedt[4]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hac0a;
    LUT4 mux_28_i6_4_lut (.A(n7[5]), .B(speedt[5]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hac0a;
    LUT4 mux_28_i7_4_lut (.A(n7[6]), .B(speedt[6]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hac0a;
    LUT4 mux_28_i8_4_lut (.A(n7[7]), .B(speedt[7]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hac0a;
    LUT4 mux_28_i9_4_lut (.A(n7[8]), .B(speedt[8]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hac0a;
    LUT4 mux_28_i10_4_lut (.A(n7[9]), .B(speedt[9]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hac0a;
    LUT4 mux_28_i11_4_lut (.A(n7[10]), .B(speedt[10]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hac0a;
    LUT4 mux_28_i12_4_lut (.A(n7[11]), .B(speedt[11]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hac0a;
    LUT4 i13779_2_lut_3_lut_4_lut (.A(stable_count[4]), .B(n21545), .C(stable_counting_N_1746), 
         .D(stable_count[5]), .Z(stable_counting_N_1759[5])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13779_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i2346_3_lut_rep_296_4_lut (.A(stable_count[4]), .B(n21545), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n21505)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2346_3_lut_rep_296_4_lut.init = 16'h7f80;
    LUT4 mux_28_i13_4_lut (.A(n7[12]), .B(speedt[12]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hac0a;
    LUT4 mux_28_i14_4_lut (.A(n7[13]), .B(speedt[13]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hac0a;
    LUT4 mux_28_i15_4_lut (.A(n7[14]), .B(speedt[14]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hac0a;
    LUT4 i14085_2_lut_rep_288_4_lut_3_lut_4_lut (.A(stable_count[4]), .B(n21545), 
         .C(stable_count[6]), .D(stable_count[5]), .Z(n21497)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i14085_2_lut_rep_288_4_lut_3_lut_4_lut.init = 16'h7ff8;
    LUT4 mux_28_i16_4_lut (.A(n7[15]), .B(speedt[15]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hac0a;
    LUT4 mux_28_i17_4_lut (.A(n7[16]), .B(speedt[16]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hac0a;
    LUT4 mux_28_i18_4_lut (.A(n7[17]), .B(speedt[17]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hac0a;
    LUT4 mux_28_i19_4_lut (.A(n7[18]), .B(speedt[18]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hac0a;
    LUT4 mux_28_i20_4_lut (.A(n7[19]), .B(speedt[19]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hac0a;
    FD1S3IX count__i1 (.D(n7[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n7[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n7[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n7[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n7[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n7[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n7[7]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n7[8]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n7[9]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n7[10]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n7[11]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n7[12]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n7[13]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n7[14]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n7[15]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n7[16]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n7[17]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n7[18]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n7[19]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX speedt__i1 (.D(n7[1]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    FD1P3IX speedt__i2 (.D(n7[2]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n7[3]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n7[4]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n7[5]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n7[6]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n7[7]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n7[8]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n7[9]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n7[10]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n7[11]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n7[12]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n7[13]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n7[14]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n7[15]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n7[16]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n7[17]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n7[18]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n7[19]), .SP(clk_1mhz_enable_66), .CD(n4298), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(hall2_old), .B(hall1_old), .C(hall2_lat), .D(hall1_lat), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(92[7:87])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i17131_3_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(stable_counting_N_1758), .Z(n19965)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i17131_3_lut.init = 16'hc8c8;
    LUT4 i2313_2_lut_rep_397 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21606)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2313_2_lut_rep_397.init = 16'h8888;
    LUT4 i2320_2_lut_rep_357_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21566)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2320_2_lut_rep_357_3_lut.init = 16'h8080;
    LUT4 i2327_2_lut_rep_336_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21545)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2327_2_lut_rep_336_3_lut_4_lut.init = 16'h8000;
    LUT4 i2325_2_lut_rep_337_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21546)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2325_2_lut_rep_337_3_lut_4_lut.init = 16'h78f0;
    LUT4 i13776_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_counting_N_1746), .D(stable_count[2]), .Z(stable_counting_N_1759[2])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13776_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i2318_2_lut_rep_358_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21567)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2318_2_lut_rep_358_3_lut.init = 16'h7878;
    LUT4 i1_2_lut_3_lut_4_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n16318)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i1_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h7ff8;
    LUT4 i13775_3_lut_rep_326 (.A(stable_count[1]), .B(stable_counting_N_1746), 
         .C(stable_count[0]), .Z(n21535)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(98[4] 103[11])
    defparam i13775_3_lut_rep_326.init = 16'h1212;
    LUT4 i5_2_lut_4_lut (.A(stable_count[1]), .B(stable_counting_N_1746), 
         .C(stable_count[0]), .D(count[19]), .Z(n17)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(98[4] 103[11])
    defparam i5_2_lut_4_lut.init = 16'h1200;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18456), 
          .S0(n7[19]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18455), .COUT(n18456), .S0(n7[17]), .S1(n7[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    LUT4 i2339_2_lut_rep_297_3_lut_4_lut (.A(stable_count[3]), .B(n21566), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21506)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2339_2_lut_rep_297_3_lut_4_lut.init = 16'h78f0;
    LUT4 i13778_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21566), .C(stable_counting_N_1746), 
         .D(stable_count[4]), .Z(stable_counting_N_1759[4])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13778_2_lut_3_lut_4_lut.init = 16'h0708;
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18454), .COUT(n18455), .S0(n7[15]), .S1(n7[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18453), .COUT(n18454), .S0(n7[13]), .S1(n7[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18452), .COUT(n18453), .S0(n7[11]), .S1(n7[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18451), .COUT(n18452), .S0(n7[9]), .S1(n7[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    LUT4 i10_4_lut (.A(n13_adj_1866), .B(n20_adj_1867), .C(count[5]), 
         .D(clk_1mhz_enable_66), .Z(n22_adj_1862)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i10_4_lut.init = 16'h8000;
    LUT4 i17167_4_lut (.A(count[13]), .B(n19989), .C(n19831), .D(count[12]), 
         .Z(n20001)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17167_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[14]), .B(stable_counting), .C(count[2]), .D(count[9]), 
         .Z(n20_adj_1867)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i17155_4_lut (.A(stable_counting_N_1759[4]), .B(n19953), .C(n13_adj_1868), 
         .D(count[0]), .Z(n19989)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17155_4_lut.init = 16'hfffe;
    LUT4 i17119_4_lut (.A(n11_adj_1869), .B(stable_counting_N_1746), .C(count[15]), 
         .D(n16318), .Z(n19953)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i17119_4_lut.init = 16'hfbfa;
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18450), 
          .COUT(n18451), .S0(n7[7]), .S1(n7[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18449), 
          .COUT(n18450), .S0(n7[5]), .S1(n7[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18448), 
          .COUT(n18449), .S0(n7[3]), .S1(n7[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18447), 
          .COUT(n18448), .S0(n7[1]), .S1(n7[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18447), 
          .S1(n7[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 mux_28_i1_4_lut (.A(n7[0]), .B(speedt[0]), .C(stable_counting_N_1758), 
         .D(n21511), .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !((C+!(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hac0a;
    LUT4 i9_4_lut (.A(n13_adj_1868), .B(n18_adj_1870), .C(count[8]), .D(count[0]), 
         .Z(n18946)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i42_2_lut (.A(count[5]), .B(count[2]), .Z(n22)) /* synthesis lut_function=(A (B)) */ ;
    defparam i42_2_lut.init = 16'h8888;
    LUT4 i8_4_lut_adj_121 (.A(n15_adj_1871), .B(n11_adj_1869), .C(count[19]), 
         .D(count[12]), .Z(n18_adj_1870)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i8_4_lut_adj_121.init = 16'hffef;
    LUT4 i5_2_lut (.A(count[15]), .B(count[13]), .Z(n15_adj_1871)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i2334_2_lut_rep_312_3_lut_4_lut (.A(stable_count[2]), .B(n21606), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21521)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2334_2_lut_rep_312_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(count[11]), .B(count[6]), .Z(n11_adj_1869)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2332_2_lut_rep_314_3_lut_4_lut (.A(stable_count[2]), .B(n21606), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21523)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2332_2_lut_rep_314_3_lut_4_lut.init = 16'h78f0;
    LUT4 i13777_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21606), .C(stable_counting_N_1746), 
         .D(stable_count[3]), .Z(stable_counting_N_1759[3])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13777_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i2_3_lut_rep_359 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_359.init = 16'hdede;
    LUT4 i3_2_lut (.A(count[7]), .B(count[10]), .Z(n13_adj_1868)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_122 (.A(count[4]), .B(count[1]), .C(count[18]), 
         .D(count[3]), .Z(n14)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_122.init = 16'h8000;
    LUT4 i17045_3_lut_4_lut (.A(count[17]), .B(count[16]), .C(count[9]), 
         .D(count[14]), .Z(n19879)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i17045_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(count[17]), .B(count[16]), .C(n14), .Z(n13_adj_1866)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    FD1S3IX count__i0 (.D(n7[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_66), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22198), .SP(stable_counting_N_1746), 
            .CD(n19965), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=302, LSE_RLINE=302 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION
//

module COMMUTATION (MB_m4_c_0, clkout_c, MC_m4_c_0, MA_m4_c_0, LED4_c, 
            enable_m4, n3175, n21589, PWM_m4, n3211, n21587, n19662, 
            n21585, free_m4, MA_m4_c_1, n3269, MC_m4_c_1, n3223, 
            MB_m4_c_1, n3187);
    output MB_m4_c_0;
    input clkout_c;
    output MC_m4_c_0;
    output MA_m4_c_0;
    output LED4_c;
    input enable_m4;
    input n3175;
    input n21589;
    input PWM_m4;
    input n3211;
    input n21587;
    input n19662;
    input n21585;
    input free_m4;
    output MA_m4_c_1;
    input n3269;
    output MC_m4_c_1;
    input n3223;
    output MB_m4_c_1;
    input n3187;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1780, n18871, n18870, n19663, clkout_c_enable_10;
    
    FD1S3IX MospairB_i1 (.D(n18871), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MB_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18870), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MC_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19663), .CK(clkout_c), .CD(led1_N_1780), 
            .Q(MA_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1P3AX led1_46 (.D(led1_N_1780), .SP(clkout_c_enable_10), .CK(clkout_c), 
            .Q(LED4_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10096_1_lut (.A(enable_m4), .Z(led1_N_1780)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i10096_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3175), .B(n21589), .C(PWM_m4), .Z(n18871)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_120 (.A(n3211), .B(n21587), .C(PWM_m4), .Z(n18870)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_120.init = 16'hbfbf;
    LUT4 i17999_3_lut (.A(n19662), .B(PWM_m4), .C(n21585), .Z(n19663)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17999_3_lut.init = 16'hbfbf;
    LUT4 i17960_2_lut (.A(free_m4), .B(enable_m4), .Z(clkout_c_enable_10)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i17960_2_lut.init = 16'h7777;
    FD1S3IX MospairA_i2 (.D(n3269), .CK(clkout_c), .CD(n19662), .Q(MA_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3211), .CK(clkout_c), .CD(n3223), .Q(MC_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3175), .CK(clkout_c), .CD(n3187), .Q(MB_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module CLKDIV
//

module CLKDIV (clk_N_683, clkout_c, clk_1mhz, pwm_clk, GND_net);
    output clk_N_683;
    input clkout_c;
    output clk_1mhz;
    output pwm_clk;
    input GND_net;
    
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(30[4:14])
    wire pi_clk /* synthesis is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(89[9:15])
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(88[9:16])
    
    wire mhz_buf, mhz_buf_N_68, pi_buf, pi_buf_N_69, pwm_buf, pwm_buf_N_67, 
        n12555, n18575;
    wire [11:0]cntpi;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(42[8:13])
    wire [8:0]n41;
    wire [4:0]count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(41[8:13])
    
    wire n19867;
    wire [4:0]n25;
    
    wire n18574, n18573, n18572, n12554, n19935, n19933, n21605;
    
    INV i18313 (.A(pi_clk), .Z(clk_N_683));
    FD1S3AX mhz_buf_29 (.D(mhz_buf_N_68), .CK(clkout_c), .Q(mhz_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(55[1] 79[8])
    defparam mhz_buf_29.GSR = "DISABLED";
    FD1S3AX pi_buf_30 (.D(pi_buf_N_69), .CK(clkout_c), .Q(pi_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(55[1] 79[8])
    defparam pi_buf_30.GSR = "DISABLED";
    FD1S3AX pwm_buf_32 (.D(pwm_buf_N_67), .CK(clkout_c), .Q(pwm_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(55[1] 79[8])
    defparam pwm_buf_32.GSR = "DISABLED";
    FD1S3AX clk_1mhz_33 (.D(mhz_buf), .CK(clkout_c), .Q(clk_1mhz)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(55[1] 79[8])
    defparam clk_1mhz_33.GSR = "DISABLED";
    FD1S3AX pwm_clk_34 (.D(pwm_buf), .CK(clkout_c), .Q(pwm_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(55[1] 79[8])
    defparam pwm_clk_34.GSR = "DISABLED";
    FD1S3AX pi_clk_35 (.D(pi_buf), .CK(clkout_c), .Q(pi_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=288, LSE_RLINE=288 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(55[1] 79[8])
    defparam pi_clk_35.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(mhz_buf), .B(n12555), .Z(mhz_buf_N_68)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    CCU2D cntpi_2060_2061_add_4_9 (.A0(cntpi[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18575), .S0(n41[7]), .S1(n41[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061_add_4_9.INIT0 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_9.INIT1 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_9.INJECT1_0 = "NO";
    defparam cntpi_2060_2061_add_4_9.INJECT1_1 = "NO";
    LUT4 i17909_4_lut (.A(count[2]), .B(count[0]), .C(count[3]), .D(n19867), 
         .Z(n12555)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(61[5:15])
    defparam i17909_4_lut.init = 16'h0400;
    LUT4 i17033_2_lut (.A(count[4]), .B(count[1]), .Z(n19867)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17033_2_lut.init = 16'h8888;
    LUT4 i15866_1_lut (.A(count[0]), .Z(n25[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam i15866_1_lut.init = 16'h5555;
    CCU2D cntpi_2060_2061_add_4_7 (.A0(cntpi[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18574), .COUT(n18575), .S0(n41[5]), .S1(n41[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061_add_4_7.INIT0 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_7.INIT1 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_7.INJECT1_0 = "NO";
    defparam cntpi_2060_2061_add_4_7.INJECT1_1 = "NO";
    CCU2D cntpi_2060_2061_add_4_5 (.A0(cntpi[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18573), .COUT(n18574), .S0(n41[3]), .S1(n41[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061_add_4_5.INIT0 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_5.INIT1 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_5.INJECT1_0 = "NO";
    defparam cntpi_2060_2061_add_4_5.INJECT1_1 = "NO";
    CCU2D cntpi_2060_2061_add_4_3 (.A0(cntpi[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18572), .COUT(n18573), .S0(n41[1]), .S1(n41[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061_add_4_3.INIT0 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_3.INIT1 = 16'hfaaa;
    defparam cntpi_2060_2061_add_4_3.INJECT1_0 = "NO";
    defparam cntpi_2060_2061_add_4_3.INJECT1_1 = "NO";
    LUT4 i15868_2_lut (.A(count[1]), .B(count[0]), .Z(n25[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam i15868_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_119 (.A(pi_buf), .B(n12554), .Z(pi_buf_N_69)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_119.init = 16'h6666;
    CCU2D cntpi_2060_2061_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18572), .S1(n41[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061_add_4_1.INIT0 = 16'hF000;
    defparam cntpi_2060_2061_add_4_1.INIT1 = 16'h0555;
    defparam cntpi_2060_2061_add_4_1.INJECT1_0 = "NO";
    defparam cntpi_2060_2061_add_4_1.INJECT1_1 = "NO";
    LUT4 i17906_4_lut (.A(n19935), .B(cntpi[2]), .C(n19933), .D(cntpi[7]), 
         .Z(n12554)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(66[5:16])
    defparam i17906_4_lut.init = 16'h0020;
    LUT4 i17101_3_lut (.A(cntpi[5]), .B(cntpi[3]), .C(cntpi[6]), .Z(n19935)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17101_3_lut.init = 16'h8080;
    LUT4 i15871_2_lut_rep_396 (.A(count[1]), .B(count[0]), .Z(n21605)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam i15871_2_lut_rep_396.init = 16'h8888;
    LUT4 i15875_2_lut_3_lut (.A(count[1]), .B(count[0]), .C(count[2]), 
         .Z(n25[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam i15875_2_lut_3_lut.init = 16'h7878;
    LUT4 i15882_2_lut_3_lut_4_lut (.A(count[1]), .B(count[0]), .C(count[3]), 
         .D(count[2]), .Z(n25[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam i15882_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i17099_4_lut (.A(cntpi[1]), .B(cntpi[0]), .C(cntpi[8]), .D(cntpi[4]), 
         .Z(n19933)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17099_4_lut.init = 16'h8000;
    LUT4 pwm_buf_I_0_1_lut (.A(pwm_buf), .Z(pwm_buf_N_67)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(73[14:25])
    defparam pwm_buf_I_0_1_lut.init = 16'h5555;
    LUT4 i15889_3_lut_4_lut (.A(count[2]), .B(n21605), .C(count[3]), .D(count[4]), 
         .Z(n25[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam i15889_3_lut_4_lut.init = 16'h7f80;
    FD1S3IX count_2059__i0 (.D(n25[0]), .CK(clkout_c), .CD(n12555), .Q(count[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam count_2059__i0.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i1 (.D(n41[0]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i1.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i2 (.D(n41[1]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i2.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i3 (.D(n41[2]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i3.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i4 (.D(n41[3]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i4.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i5 (.D(n41[4]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i5.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i6 (.D(n41[5]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i6.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i7 (.D(n41[6]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i7.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i8 (.D(n41[7]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i8.GSR = "DISABLED";
    FD1S3IX cntpi_2060_2061__i9 (.D(n41[8]), .CK(clkout_c), .CD(n12554), 
            .Q(cntpi[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(57[11:16])
    defparam cntpi_2060_2061__i9.GSR = "DISABLED";
    FD1S3IX count_2059__i1 (.D(n25[1]), .CK(clkout_c), .CD(n12555), .Q(count[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam count_2059__i1.GSR = "DISABLED";
    FD1S3IX count_2059__i2 (.D(n25[2]), .CK(clkout_c), .CD(n12555), .Q(count[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam count_2059__i2.GSR = "DISABLED";
    FD1S3IX count_2059__i3 (.D(n25[3]), .CK(clkout_c), .CD(n12555), .Q(count[3]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam count_2059__i3.GSR = "DISABLED";
    FD1S3IX count_2059__i4 (.D(n25[4]), .CK(clkout_c), .CD(n12555), .Q(count[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/clockdivider.vhd(56[11:16])
    defparam count_2059__i4.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U0
//

module PWMGENERATOR_U0 (PWM_m3, pwm_clk, free_m3, clkout_c_enable_176, 
            hallsense_m3, n21591, enable_m3, n3093, PWMdut_m3, GND_net, 
            n21592, n19650, n21593, n3057);
    output PWM_m3;
    input pwm_clk;
    output free_m3;
    input clkout_c_enable_176;
    input [2:0]hallsense_m3;
    output n21591;
    input enable_m3;
    output n3093;
    input [9:0]PWMdut_m3;
    input GND_net;
    output n21592;
    output n19650;
    output n21593;
    output n3057;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_1805, free_N_1817, n17;
    wire [9:0]cnt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(41[10:13])
    
    wire n16, n12551, n18526, n3674, n18525, n7, n18524, n18523, 
        n9, n10, n18522, n18546;
    wire [9:0]n45;
    
    wire n18545, n18544, n18543, n18542, n10_adj_1860, n10961, n14, 
        n10_adj_1861;
    
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m3)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=328, LSE_RLINE=328 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_176), .CK(pwm_clk), 
            .Q(free_m3));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i17897_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n12551)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(73[6:16])
    defparam i17897_4_lut.init = 16'h0400;
    LUT4 i1629_3_lut_rep_382 (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .Z(n21591)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1629_3_lut_rep_382.init = 16'h1414;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i17941_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .D(enable_m3), .Z(n3093)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17941_2_lut_4_lut.init = 16'hebff;
    LUT4 i6_4_lut (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut.init = 16'hffef;
    CCU2D sub_1793_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m3[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18526), .S1(n3674));
    defparam sub_1793_add_2_11.INIT0 = 16'h5999;
    defparam sub_1793_add_2_11.INIT1 = 16'h0000;
    defparam sub_1793_add_2_11.INJECT1_0 = "NO";
    defparam sub_1793_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1793_add_2_9 (.A0(PWMdut_m3[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m3[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18525), 
          .COUT(n18526));
    defparam sub_1793_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1793_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1793_add_2_9.INJECT1_0 = "NO";
    defparam sub_1793_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1793_add_2_7 (.A0(PWMdut_m3[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m3[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18524), 
          .COUT(n18525));
    defparam sub_1793_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1793_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1793_add_2_7.INJECT1_0 = "NO";
    defparam sub_1793_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1793_add_2_5 (.A0(PWMdut_m3[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m3[4]), .C1(n9), .D1(n10), .CIN(n18523), 
          .COUT(n18524));
    defparam sub_1793_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1793_add_2_5.INIT1 = 16'h5999;
    defparam sub_1793_add_2_5.INJECT1_0 = "NO";
    defparam sub_1793_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_383 (.A(enable_m3), .B(free_m3), .Z(n21592)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1_2_lut_rep_383.init = 16'h2222;
    LUT4 i17945_3_lut_4_lut (.A(enable_m3), .B(free_m3), .C(hallsense_m3[2]), 
         .D(hallsense_m3[0]), .Z(n19650)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17945_3_lut_4_lut.init = 16'hfddf;
    LUT4 i1599_3_lut_rep_384 (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .Z(n21593)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1599_3_lut_rep_384.init = 16'h1414;
    LUT4 i17938_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .D(enable_m3), .Z(n3057)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17938_2_lut_4_lut.init = 16'hebff;
    CCU2D sub_1793_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m3[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m3[2]), .C1(n9), .D1(n10), .CIN(n18522), 
          .COUT(n18523));
    defparam sub_1793_add_2_3.INIT0 = 16'h5999;
    defparam sub_1793_add_2_3.INIT1 = 16'h5999;
    defparam sub_1793_add_2_3.INJECT1_0 = "NO";
    defparam sub_1793_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1793_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m3[0]), .C1(n9), .D1(n10), 
          .COUT(n18522));
    defparam sub_1793_add_2_1.INIT0 = 16'h0000;
    defparam sub_1793_add_2_1.INIT1 = 16'h5999;
    defparam sub_1793_add_2_1.INJECT1_0 = "NO";
    defparam sub_1793_add_2_1.INJECT1_1 = "NO";
    CCU2D cnt_2066_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18546), .S0(n45[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2066_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2066_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18545), 
          .COUT(n18546), .S0(n45[7]), .S1(n45[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2066_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18544), 
          .COUT(n18545), .S0(n45[5]), .S1(n45[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2066_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18543), 
          .COUT(n18544), .S0(n45[3]), .S1(n45[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2066_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18542), 
          .COUT(n18543), .S0(n45[1]), .S1(n45[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2066_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2066_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_3.INJECT1_1 = "NO";
    LUT4 i2_3_lut (.A(PWMdut_m3[5]), .B(PWMdut_m3[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_1860), .B(PWMdut_m3[9]), .C(PWMdut_m3[8]), 
         .D(PWMdut_m3[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2259_3_lut (.A(n10961), .B(PWMdut_m3[4]), .C(PWMdut_m3[3]), 
         .Z(n10_adj_1860)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2259_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D cnt_2066_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18542), .S1(n45[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2066_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2066_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2066_add_4_1.INJECT1_1 = "NO";
    LUT4 i1795_1_lut (.A(n3674), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1795_1_lut.init = 16'h5555;
    LUT4 i17877_4_lut (.A(PWMdut_m3[5]), .B(n14), .C(n10_adj_1861), .D(PWMdut_m3[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i17877_4_lut.init = 16'h0001;
    LUT4 i6_4_lut_adj_117 (.A(PWMdut_m3[9]), .B(PWMdut_m3[3]), .C(PWMdut_m3[4]), 
         .D(n10961), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut_adj_117.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[7]), .Z(n10_adj_1861)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_118 (.A(PWMdut_m3[2]), .B(PWMdut_m3[1]), .C(PWMdut_m3[0]), 
         .Z(n10961)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_118.init = 16'hfefe;
    FD1S3IX cnt_2066__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12551), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i0.GSR = "ENABLED";
    FD1S3IX cnt_2066__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12551), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i1.GSR = "ENABLED";
    FD1S3IX cnt_2066__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12551), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i2.GSR = "ENABLED";
    FD1S3IX cnt_2066__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12551), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i3.GSR = "ENABLED";
    FD1S3IX cnt_2066__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12551), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i4.GSR = "ENABLED";
    FD1S3IX cnt_2066__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12551), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i5.GSR = "ENABLED";
    FD1S3IX cnt_2066__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12551), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i6.GSR = "ENABLED";
    FD1S3IX cnt_2066__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12551), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i7.GSR = "ENABLED";
    FD1S3IX cnt_2066__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12551), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i8.GSR = "ENABLED";
    FD1S3IX cnt_2066__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12551), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2066__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U1
//

module PWMGENERATOR_U1 (PWM_m2, pwm_clk, free_m2, clkout_c_enable_176, 
            PWMdut_m2, GND_net, hallsense_m2, n21596, enable_m2, n2963, 
            n21598, n2927);
    output PWM_m2;
    input pwm_clk;
    output free_m2;
    input clkout_c_enable_176;
    input [9:0]PWMdut_m2;
    input GND_net;
    input [2:0]hallsense_m2;
    output n21596;
    input enable_m2;
    output n2963;
    output n21598;
    output n2927;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_1805, free_N_1817, n18531;
    wire [9:0]cnt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(41[10:13])
    
    wire n3661, n18530, n7, n19981, n6, n12552, n19937, n18529, 
        n18528, n9, n10, n18527, n10_adj_1858, n10965, n18551;
    wire [9:0]n45;
    
    wire n18550, n18549, n18548, n18547, n14, n10_adj_1859;
    
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m2)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=318, LSE_RLINE=318 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_176), .CK(pwm_clk), 
            .Q(free_m2));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    CCU2D sub_1791_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m2[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18531), .S1(n3661));
    defparam sub_1791_add_2_11.INIT0 = 16'h5999;
    defparam sub_1791_add_2_11.INIT1 = 16'h0000;
    defparam sub_1791_add_2_11.INJECT1_0 = "NO";
    defparam sub_1791_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1791_add_2_9 (.A0(PWMdut_m2[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m2[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18530), 
          .COUT(n18531));
    defparam sub_1791_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1791_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1791_add_2_9.INJECT1_0 = "NO";
    defparam sub_1791_add_2_9.INJECT1_1 = "NO";
    LUT4 i17900_4_lut (.A(cnt[0]), .B(n19981), .C(cnt[2]), .D(n6), .Z(n12552)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(73[6:16])
    defparam i17900_4_lut.init = 16'h0004;
    LUT4 i17147_3_lut (.A(cnt[7]), .B(n19937), .C(cnt[3]), .Z(n19981)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17147_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i17103_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n19937)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17103_4_lut.init = 16'h8000;
    CCU2D sub_1791_add_2_7 (.A0(PWMdut_m2[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m2[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18529), 
          .COUT(n18530));
    defparam sub_1791_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1791_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1791_add_2_7.INJECT1_0 = "NO";
    defparam sub_1791_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1791_add_2_5 (.A0(PWMdut_m2[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m2[4]), .C1(n9), .D1(n10), .CIN(n18528), 
          .COUT(n18529));
    defparam sub_1791_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1791_add_2_5.INIT1 = 16'h5999;
    defparam sub_1791_add_2_5.INJECT1_0 = "NO";
    defparam sub_1791_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1791_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m2[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m2[2]), .C1(n9), .D1(n10), .CIN(n18527), 
          .COUT(n18528));
    defparam sub_1791_add_2_3.INIT0 = 16'h5999;
    defparam sub_1791_add_2_3.INIT1 = 16'h5999;
    defparam sub_1791_add_2_3.INJECT1_0 = "NO";
    defparam sub_1791_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1791_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m2[0]), .C1(n9), .D1(n10), 
          .COUT(n18527));
    defparam sub_1791_add_2_1.INIT0 = 16'h0000;
    defparam sub_1791_add_2_1.INIT1 = 16'h5999;
    defparam sub_1791_add_2_1.INJECT1_0 = "NO";
    defparam sub_1791_add_2_1.INJECT1_1 = "NO";
    LUT4 i1537_3_lut_rep_387 (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .Z(n21596)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1537_3_lut_rep_387.init = 16'h1414;
    LUT4 i17931_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .D(enable_m2), .Z(n2963)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17931_2_lut_4_lut.init = 16'hebff;
    LUT4 i2_3_lut (.A(PWMdut_m2[5]), .B(PWMdut_m2[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_1858), .B(PWMdut_m2[9]), .C(PWMdut_m2[8]), 
         .D(PWMdut_m2[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2262_3_lut (.A(n10965), .B(PWMdut_m2[4]), .C(PWMdut_m2[3]), 
         .Z(n10_adj_1858)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2262_3_lut.init = 16'hecec;
    LUT4 i1507_3_lut_rep_389 (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .Z(n21598)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1507_3_lut_rep_389.init = 16'h1414;
    LUT4 i17928_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .D(enable_m2), .Z(n2927)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17928_2_lut_4_lut.init = 16'hebff;
    CCU2D cnt_2065_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18551), .S0(n45[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2065_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18550), 
          .COUT(n18551), .S0(n45[7]), .S1(n45[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18549), 
          .COUT(n18550), .S0(n45[5]), .S1(n45[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18548), 
          .COUT(n18549), .S0(n45[3]), .S1(n45[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18547), 
          .COUT(n18548), .S0(n45[1]), .S1(n45[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2065_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2065_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2065_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18547), .S1(n45[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2065_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2065_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2065_add_4_1.INJECT1_1 = "NO";
    LUT4 i3_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1793_1_lut (.A(n3661), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1793_1_lut.init = 16'h5555;
    LUT4 i17832_4_lut (.A(PWMdut_m2[5]), .B(n14), .C(n10_adj_1859), .D(PWMdut_m2[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i17832_4_lut.init = 16'h0001;
    FD1S3IX cnt_2065__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12552), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i0.GSR = "ENABLED";
    LUT4 i6_4_lut (.A(PWMdut_m2[9]), .B(PWMdut_m2[3]), .C(PWMdut_m2[4]), 
         .D(n10965), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[7]), .Z(n10_adj_1859)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_116 (.A(PWMdut_m2[2]), .B(PWMdut_m2[1]), .C(PWMdut_m2[0]), 
         .Z(n10965)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_116.init = 16'hfefe;
    FD1S3IX cnt_2065__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12552), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i1.GSR = "ENABLED";
    FD1S3IX cnt_2065__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12552), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i2.GSR = "ENABLED";
    FD1S3IX cnt_2065__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12552), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i3.GSR = "ENABLED";
    FD1S3IX cnt_2065__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12552), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i4.GSR = "ENABLED";
    FD1S3IX cnt_2065__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12552), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i5.GSR = "ENABLED";
    FD1S3IX cnt_2065__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12552), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i6.GSR = "ENABLED";
    FD1S3IX cnt_2065__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12552), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i7.GSR = "ENABLED";
    FD1S3IX cnt_2065__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12552), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i8.GSR = "ENABLED";
    FD1S3IX cnt_2065__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12552), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2065__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U2
//

module PWMGENERATOR_U2 (GND_net, PWMdut_m1, PWM_m1, pwm_clk, free_m1, 
            clkout_c_enable_164, hallsense_m1, n21573, enable_m1, n2833, 
            n21574, n19654, n21575, n2797);
    input GND_net;
    input [9:0]PWMdut_m1;
    output PWM_m1;
    input pwm_clk;
    output free_m1;
    input clkout_c_enable_164;
    input [2:0]hallsense_m1;
    output n21573;
    input enable_m1;
    output n2833;
    output n21574;
    output n19654;
    output n21575;
    output n2797;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(88[9:16])
    wire [9:0]cnt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(41[10:13])
    
    wire n9, n10, n18532, PWM_N_1805, free_N_1817, n7, n19995, 
        n6, n12553, n19971, n18556;
    wire [9:0]n45;
    
    wire n18555, n18554, n18553, n18552, n10_adj_1856, n10963, n14, 
        n10_adj_1857, n18536, n3648, n18535, n18534, n18533;
    
    CCU2D sub_1789_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m1[0]), .C1(n9), .D1(n10), 
          .COUT(n18532));
    defparam sub_1789_add_2_1.INIT0 = 16'h0000;
    defparam sub_1789_add_2_1.INIT1 = 16'h5999;
    defparam sub_1789_add_2_1.INJECT1_0 = "NO";
    defparam sub_1789_add_2_1.INJECT1_1 = "NO";
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=308, LSE_RLINE=308 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_164), .CK(pwm_clk), 
            .Q(free_m1));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(PWMdut_m1[5]), .B(PWMdut_m1[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i17903_4_lut (.A(cnt[0]), .B(n19995), .C(cnt[2]), .D(n6), .Z(n12553)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(73[6:16])
    defparam i17903_4_lut.init = 16'h0004;
    LUT4 i17161_3_lut (.A(cnt[7]), .B(n19971), .C(cnt[3]), .Z(n19995)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17161_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i17137_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n19971)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17137_4_lut.init = 16'h8000;
    CCU2D cnt_2064_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18556), .S0(n45[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2064_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2064_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2064_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2064_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18555), 
          .COUT(n18556), .S0(n45[7]), .S1(n45[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2064_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2064_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2064_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2064_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18554), 
          .COUT(n18555), .S0(n45[5]), .S1(n45[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2064_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2064_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2064_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2064_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18553), 
          .COUT(n18554), .S0(n45[3]), .S1(n45[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2064_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2064_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2064_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2064_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18552), 
          .COUT(n18553), .S0(n45[1]), .S1(n45[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2064_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2064_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2064_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2064_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18552), .S1(n45[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2064_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2064_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2064_add_4_1.INJECT1_1 = "NO";
    LUT4 i3_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i3_4_lut (.A(n10_adj_1856), .B(PWMdut_m1[9]), .C(PWMdut_m1[8]), 
         .D(PWMdut_m1[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2265_3_lut (.A(n10963), .B(PWMdut_m1[4]), .C(PWMdut_m1[3]), 
         .Z(n10_adj_1856)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2265_3_lut.init = 16'hecec;
    LUT4 i2_3_lut_adj_115 (.A(PWMdut_m1[2]), .B(PWMdut_m1[1]), .C(PWMdut_m1[0]), 
         .Z(n10963)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_115.init = 16'hfefe;
    LUT4 i17835_4_lut (.A(PWMdut_m1[5]), .B(n14), .C(n10_adj_1857), .D(PWMdut_m1[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i17835_4_lut.init = 16'h0001;
    CCU2D sub_1789_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m1[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18536), .S1(n3648));
    defparam sub_1789_add_2_11.INIT0 = 16'h5999;
    defparam sub_1789_add_2_11.INIT1 = 16'h0000;
    defparam sub_1789_add_2_11.INJECT1_0 = "NO";
    defparam sub_1789_add_2_11.INJECT1_1 = "NO";
    LUT4 i6_4_lut (.A(PWMdut_m1[9]), .B(PWMdut_m1[3]), .C(PWMdut_m1[4]), 
         .D(n10963), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    CCU2D sub_1789_add_2_9 (.A0(PWMdut_m1[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m1[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18535), 
          .COUT(n18536));
    defparam sub_1789_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1789_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1789_add_2_9.INJECT1_0 = "NO";
    defparam sub_1789_add_2_9.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[7]), .Z(n10_adj_1857)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    CCU2D sub_1789_add_2_7 (.A0(PWMdut_m1[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m1[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18534), 
          .COUT(n18535));
    defparam sub_1789_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1789_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1789_add_2_7.INJECT1_0 = "NO";
    defparam sub_1789_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1789_add_2_5 (.A0(PWMdut_m1[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m1[4]), .C1(n9), .D1(n10), .CIN(n18533), 
          .COUT(n18534));
    defparam sub_1789_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1789_add_2_5.INIT1 = 16'h5999;
    defparam sub_1789_add_2_5.INJECT1_0 = "NO";
    defparam sub_1789_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1789_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m1[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m1[2]), .C1(n9), .D1(n10), .CIN(n18532), 
          .COUT(n18533));
    defparam sub_1789_add_2_3.INIT0 = 16'h5999;
    defparam sub_1789_add_2_3.INIT1 = 16'h5999;
    defparam sub_1789_add_2_3.INJECT1_0 = "NO";
    defparam sub_1789_add_2_3.INJECT1_1 = "NO";
    LUT4 i1445_3_lut_rep_364 (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .Z(n21573)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1445_3_lut_rep_364.init = 16'h1414;
    LUT4 i17921_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .D(enable_m1), .Z(n2833)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17921_2_lut_4_lut.init = 16'hebff;
    LUT4 i1_2_lut_rep_365 (.A(enable_m1), .B(free_m1), .Z(n21574)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1_2_lut_rep_365.init = 16'h2222;
    LUT4 i17925_3_lut_4_lut (.A(enable_m1), .B(free_m1), .C(hallsense_m1[2]), 
         .D(hallsense_m1[0]), .Z(n19654)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17925_3_lut_4_lut.init = 16'hfddf;
    LUT4 i1415_3_lut_rep_366 (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .Z(n21575)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1415_3_lut_rep_366.init = 16'h1414;
    LUT4 i17918_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .D(enable_m1), .Z(n2797)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17918_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2064__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12553), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i0.GSR = "ENABLED";
    LUT4 i1791_1_lut (.A(n3648), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1791_1_lut.init = 16'h5555;
    FD1S3IX cnt_2064__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12553), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i1.GSR = "ENABLED";
    FD1S3IX cnt_2064__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12553), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i2.GSR = "ENABLED";
    FD1S3IX cnt_2064__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12553), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i3.GSR = "ENABLED";
    FD1S3IX cnt_2064__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12553), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i4.GSR = "ENABLED";
    FD1S3IX cnt_2064__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12553), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i5.GSR = "ENABLED";
    FD1S3IX cnt_2064__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12553), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i6.GSR = "ENABLED";
    FD1S3IX cnt_2064__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12553), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i7.GSR = "ENABLED";
    FD1S3IX cnt_2064__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12553), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i8.GSR = "ENABLED";
    FD1S3IX cnt_2064__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12553), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2064__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \PID(16000000,160000000,10000000) 
//

module \PID(16000000,160000000,10000000)  (clk_N_683, GND_net, PWMdut_m3, 
            dir_m2, dir_m3, dir_m1, dir_m4, speed_set_m2, speed_set_m1, 
            VCC_net, speed_set_m4, \speed_m4[0] , \speed_m3[0] , n21544, 
            n4132, \speed_m3[3] , \speed_m2[3] , \speed_m4[12] , \speed_m3[7] , 
            \speed_m2[7] , \speed_m3[8] , \speed_m2[8] , \speed_m3[9] , 
            \speed_m2[9] , \speed_m3[12] , \speed_m2[12] , \speed_m4[9] , 
            \speed_m4[8] , \speed_m4[18] , \speed_m3[18] , \speed_m4[7] , 
            \speed_m4[3] , \speed_m4[17] , \speed_m3[17] , \speed_m4[16] , 
            \speed_m3[16] , \speed_m4[15] , \speed_m3[15] , \speed_m4[14] , 
            \speed_m3[14] , \speed_m4[13] , \speed_m3[13] , \speed_m4[11] , 
            \speed_m3[11] , \speed_m4[10] , \speed_m3[10] , \speed_m4[6] , 
            \speed_m3[6] , \speed_m4[5] , \speed_m3[5] , \speed_m4[4] , 
            \speed_m3[4] , \speed_m4[2] , \speed_m3[2] , n22203, \speed_m4[1] , 
            \speed_m3[1] , \speed_m1[0] , \speed_m2[0] , \speed_m1[18] , 
            \speed_m2[18] , \speed_m1[17] , \speed_m2[17] , \speed_m1[16] , 
            \speed_m2[16] , \speed_m1[15] , \speed_m2[15] , \speed_m1[14] , 
            \speed_m2[14] , \speed_m1[13] , \speed_m2[13] , \speed_m1[11] , 
            \speed_m2[11] , \speed_m1[10] , \speed_m2[10] , \speed_m1[6] , 
            \speed_m2[6] , \speed_m1[5] , \speed_m2[5] , \speed_m1[4] , 
            \speed_m2[4] , \speed_m1[2] , \speed_m2[2] , \speed_m1[1] , 
            \speed_m2[1] , \speed_m1[19] , \speed_m2[19] , n5, \speed_m1[12] , 
            \speed_m1[9] , \speed_m1[8] , \speed_m1[7] , \speed_m1[3] , 
            PWMdut_m2, PWMdut_m1, speed_set_m3, n7, n20183, PWMdut_m4);
    input clk_N_683;
    input GND_net;
    output [9:0]PWMdut_m3;
    output dir_m2;
    output dir_m3;
    output dir_m1;
    output dir_m4;
    input [20:0]speed_set_m2;
    input [20:0]speed_set_m1;
    input VCC_net;
    input [20:0]speed_set_m4;
    input \speed_m4[0] ;
    input \speed_m3[0] ;
    output n21544;
    output n4132;
    input \speed_m3[3] ;
    input \speed_m2[3] ;
    input \speed_m4[12] ;
    input \speed_m3[7] ;
    input \speed_m2[7] ;
    input \speed_m3[8] ;
    input \speed_m2[8] ;
    input \speed_m3[9] ;
    input \speed_m2[9] ;
    input \speed_m3[12] ;
    input \speed_m2[12] ;
    input \speed_m4[9] ;
    input \speed_m4[8] ;
    input \speed_m4[18] ;
    input \speed_m3[18] ;
    input \speed_m4[7] ;
    input \speed_m4[3] ;
    input \speed_m4[17] ;
    input \speed_m3[17] ;
    input \speed_m4[16] ;
    input \speed_m3[16] ;
    input \speed_m4[15] ;
    input \speed_m3[15] ;
    input \speed_m4[14] ;
    input \speed_m3[14] ;
    input \speed_m4[13] ;
    input \speed_m3[13] ;
    input \speed_m4[11] ;
    input \speed_m3[11] ;
    input \speed_m4[10] ;
    input \speed_m3[10] ;
    input \speed_m4[6] ;
    input \speed_m3[6] ;
    input \speed_m4[5] ;
    input \speed_m3[5] ;
    input \speed_m4[4] ;
    input \speed_m3[4] ;
    input \speed_m4[2] ;
    input \speed_m3[2] ;
    input n22203;
    input \speed_m4[1] ;
    input \speed_m3[1] ;
    input \speed_m1[0] ;
    input \speed_m2[0] ;
    input \speed_m1[18] ;
    input \speed_m2[18] ;
    input \speed_m1[17] ;
    input \speed_m2[17] ;
    input \speed_m1[16] ;
    input \speed_m2[16] ;
    input \speed_m1[15] ;
    input \speed_m2[15] ;
    input \speed_m1[14] ;
    input \speed_m2[14] ;
    input \speed_m1[13] ;
    input \speed_m2[13] ;
    input \speed_m1[11] ;
    input \speed_m2[11] ;
    input \speed_m1[10] ;
    input \speed_m2[10] ;
    input \speed_m1[6] ;
    input \speed_m2[6] ;
    input \speed_m1[5] ;
    input \speed_m2[5] ;
    input \speed_m1[4] ;
    input \speed_m2[4] ;
    input \speed_m1[2] ;
    input \speed_m2[2] ;
    input \speed_m1[1] ;
    input \speed_m2[1] ;
    input \speed_m1[19] ;
    input \speed_m2[19] ;
    output n5;
    input \speed_m1[12] ;
    input \speed_m1[9] ;
    input \speed_m1[8] ;
    input \speed_m1[7] ;
    input \speed_m1[3] ;
    output [9:0]PWMdut_m2;
    output [9:0]PWMdut_m1;
    input [20:0]speed_set_m3;
    input n7;
    output n20183;
    output [9:0]PWMdut_m4;
    
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(30[4:14])
    wire [28:0]backOut0;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(77[9:17])
    
    wire clk_N_683_enable_73;
    wire [28:0]backOut1_28__N_1445;
    wire [28:0]backOut1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(78[9:17])
    
    wire clk_N_683_enable_41;
    wire [28:0]multOut;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(88[9:16])
    wire [53:0]multOut_28__N_1178;
    wire [28:0]intgOut0;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(67[9:17])
    
    wire clk_N_683_enable_101;
    wire [28:0]intgOut1_28__N_766;
    wire [28:0]intgOut1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(68[9:17])
    
    wire clk_N_683_enable_129;
    wire [28:0]intgOut2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(69[9:17])
    
    wire clk_N_683_enable_157;
    wire [28:0]intgOut3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(70[9:17])
    
    wire clk_N_683_enable_185;
    wire [28:0]Out0;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(72[9:13])
    
    wire clk_N_683_enable_213;
    wire [28:0]Out1;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(73[9:13])
    
    wire clk_N_683_enable_241;
    wire [28:0]Out2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(74[9:13])
    
    wire clk_N_683_enable_269;
    wire [28:0]Out3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(75[9:13])
    
    wire clk_N_683_enable_297;
    wire [28:0]backOut2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(79[9:17])
    
    wire clk_N_683_enable_325;
    wire [28:0]backOut3;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(80[9:17])
    
    wire clk_N_683_enable_353, n18711;
    wire [28:0]addOut;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(92[9:15])
    
    wire n18712;
    wire [24:0]subOut;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(84[9:15])
    wire [25:0]subOut_24__N_1135;
    
    wire n18710;
    wire [28:0]backOut0_28__N_1416;
    wire [28:0]backOut2_28__N_1474;
    
    wire clk_N_683_enable_392, n12655;
    wire [9:0]n2176;
    wire [4:0]ss;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(96[9:11])
    
    wire n14, n15, n19725, n21572, n21571, n18412, n5171, n5173;
    wire [21:0]n2244;
    
    wire n18413, subIn1_24__N_1300, dirout_m3_N_1578, subIn1_24__N_1113, 
        dirout_m4_N_1581, n21554, n21549, n20450, n21550, n21578, 
        n21522, n22208, n21613, n21612, n4138, n20179, n5129, 
        n5087, n2436, n5177, n35, n21500, n5704, n920, n3635;
    wire [28:0]intgOut0_28__N_735;
    
    wire n5690, n5692, n5694;
    wire [28:0]n648;
    
    wire n21551;
    wire [28:0]n678;
    
    wire n21524, n15859;
    wire [28:0]n558;
    
    wire n5127, n5085, n5175, n5696, n5698, n5706, n5708, n5125, 
        n5083, n5123, n5081, n14_adj_1826, n10, n18862, n5710, 
        n5712, n6, n18863, n5121, n5079, n5169, n5728, n5714, 
        n5253, n5119, n5077, n5167, n5688, n5720, n5702, n5700, 
        n5716, n5718, n5722, n5117, n5075, n5165, n22196, n22199, 
        n42, n21499, n21484, n5724, n18709, n21483, n5115, n5073, 
        n5163, n5113, n5071, n5161, n18708, n14_adj_1827, n10_adj_1828, 
        n18821, n5111, n5069, n5159, n6_adj_1829, n18822;
    wire [23:0]multIn2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(87[9:16])
    
    wire mult_29s_25s_0_pp_1_2, mult_29s_25s_0_pp_2_4, mult_29s_25s_0_pp_3_6, 
        mult_29s_25s_0_pp_4_8, mult_29s_25s_0_pp_5_10, mult_29s_25s_0_pp_6_12, 
        mult_29s_25s_0_pp_7_14, mult_29s_25s_0_pp_8_16, mult_29s_25s_0_pp_9_18, 
        mult_29s_25s_0_pp_10_20, mult_29s_25s_0_pp_11_22, mult_29s_25s_0_pp_12_24, 
        mult_29s_25s_0_pp_12_25, mult_29s_25s_0_pp_12_26, mult_29s_25s_0_pp_12_27, 
        mult_29s_25s_0_pp_12_28, mult_29s_25s_0_cin_lr_2, mult_29s_25s_0_cin_lr_4, 
        mult_29s_25s_0_cin_lr_6, mult_29s_25s_0_cin_lr_8, mult_29s_25s_0_cin_lr_10, 
        mult_29s_25s_0_cin_lr_12, mult_29s_25s_0_cin_lr_14, mult_29s_25s_0_cin_lr_16, 
        mult_29s_25s_0_cin_lr_18, mult_29s_25s_0_cin_lr_20, mult_29s_25s_0_cin_lr_22, 
        co_mult_29s_25s_0_0_1, mult_29s_25s_0_pp_0_2, co_mult_29s_25s_0_0_2, 
        s_mult_29s_25s_0_0_4, mult_29s_25s_0_pp_0_4, mult_29s_25s_0_pp_0_3, 
        mult_29s_25s_0_pp_1_4, mult_29s_25s_0_pp_1_3, co_mult_29s_25s_0_0_3, 
        s_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_6, mult_29s_25s_0_pp_0_6, 
        mult_29s_25s_0_pp_0_5, mult_29s_25s_0_pp_1_6, mult_29s_25s_0_pp_1_5, 
        co_mult_29s_25s_0_0_4, s_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_8, 
        mult_29s_25s_0_pp_0_8, mult_29s_25s_0_pp_0_7, mult_29s_25s_0_pp_1_8, 
        mult_29s_25s_0_pp_1_7, co_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_10, mult_29s_25s_0_pp_0_10, mult_29s_25s_0_pp_0_9, 
        mult_29s_25s_0_pp_1_10, mult_29s_25s_0_pp_1_9, co_mult_29s_25s_0_0_6, 
        s_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_12, mult_29s_25s_0_pp_0_12, 
        mult_29s_25s_0_pp_0_11, mult_29s_25s_0_pp_1_12, mult_29s_25s_0_pp_1_11, 
        co_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_14, 
        mult_29s_25s_0_pp_0_14, mult_29s_25s_0_pp_0_13, mult_29s_25s_0_pp_1_14, 
        mult_29s_25s_0_pp_1_13, co_mult_29s_25s_0_0_8, s_mult_29s_25s_0_0_15, 
        s_mult_29s_25s_0_0_16, mult_29s_25s_0_pp_0_16, mult_29s_25s_0_pp_0_15, 
        mult_29s_25s_0_pp_1_16, mult_29s_25s_0_pp_1_15, co_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_17, s_mult_29s_25s_0_0_18, mult_29s_25s_0_pp_0_18, 
        mult_29s_25s_0_pp_0_17, mult_29s_25s_0_pp_1_18, mult_29s_25s_0_pp_1_17, 
        co_mult_29s_25s_0_0_10, s_mult_29s_25s_0_0_19, s_mult_29s_25s_0_0_20, 
        mult_29s_25s_0_pp_0_20, mult_29s_25s_0_pp_0_19, mult_29s_25s_0_pp_1_20, 
        mult_29s_25s_0_pp_1_19, co_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_21, 
        s_mult_29s_25s_0_0_22, mult_29s_25s_0_pp_0_22, mult_29s_25s_0_pp_0_21, 
        mult_29s_25s_0_pp_1_22, mult_29s_25s_0_pp_1_21, co_mult_29s_25s_0_0_12, 
        s_mult_29s_25s_0_0_23, s_mult_29s_25s_0_0_24, mult_29s_25s_0_pp_0_24, 
        mult_29s_25s_0_pp_0_23, mult_29s_25s_0_pp_1_24, mult_29s_25s_0_pp_1_23, 
        co_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_25, s_mult_29s_25s_0_0_26, 
        mult_29s_25s_0_pp_0_26, mult_29s_25s_0_pp_0_25, mult_29s_25s_0_pp_1_26, 
        mult_29s_25s_0_pp_1_25, s_mult_29s_25s_0_0_27, s_mult_29s_25s_0_0_28, 
        mult_29s_25s_0_pp_0_28, mult_29s_25s_0_pp_0_27, mult_29s_25s_0_pp_1_28, 
        mult_29s_25s_0_pp_1_27, co_mult_29s_25s_0_1_1, s_mult_29s_25s_0_1_6, 
        mult_29s_25s_0_pp_2_6, co_mult_29s_25s_0_1_2, s_mult_29s_25s_0_1_7, 
        s_mult_29s_25s_0_1_8, mult_29s_25s_0_pp_2_8, mult_29s_25s_0_pp_2_7, 
        mult_29s_25s_0_pp_3_8, mult_29s_25s_0_pp_3_7, co_mult_29s_25s_0_1_3, 
        s_mult_29s_25s_0_1_9, s_mult_29s_25s_0_1_10, mult_29s_25s_0_pp_2_10, 
        mult_29s_25s_0_pp_2_9, mult_29s_25s_0_pp_3_10, mult_29s_25s_0_pp_3_9, 
        co_mult_29s_25s_0_1_4, s_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_12, 
        mult_29s_25s_0_pp_2_12, mult_29s_25s_0_pp_2_11, mult_29s_25s_0_pp_3_12, 
        mult_29s_25s_0_pp_3_11, co_mult_29s_25s_0_1_5, s_mult_29s_25s_0_1_13, 
        s_mult_29s_25s_0_1_14, mult_29s_25s_0_pp_2_14, mult_29s_25s_0_pp_2_13, 
        mult_29s_25s_0_pp_3_14, mult_29s_25s_0_pp_3_13, co_mult_29s_25s_0_1_6, 
        s_mult_29s_25s_0_1_15, s_mult_29s_25s_0_1_16, mult_29s_25s_0_pp_2_16, 
        mult_29s_25s_0_pp_2_15, mult_29s_25s_0_pp_3_16, mult_29s_25s_0_pp_3_15, 
        co_mult_29s_25s_0_1_7, s_mult_29s_25s_0_1_17, s_mult_29s_25s_0_1_18, 
        mult_29s_25s_0_pp_2_18, mult_29s_25s_0_pp_2_17, mult_29s_25s_0_pp_3_18, 
        mult_29s_25s_0_pp_3_17, co_mult_29s_25s_0_1_8, s_mult_29s_25s_0_1_19, 
        s_mult_29s_25s_0_1_20, mult_29s_25s_0_pp_2_20, mult_29s_25s_0_pp_2_19, 
        mult_29s_25s_0_pp_3_20, mult_29s_25s_0_pp_3_19, co_mult_29s_25s_0_1_9, 
        s_mult_29s_25s_0_1_21, s_mult_29s_25s_0_1_22, mult_29s_25s_0_pp_2_22, 
        mult_29s_25s_0_pp_2_21, mult_29s_25s_0_pp_3_22, mult_29s_25s_0_pp_3_21, 
        co_mult_29s_25s_0_1_10, s_mult_29s_25s_0_1_23, s_mult_29s_25s_0_1_24, 
        mult_29s_25s_0_pp_2_24, mult_29s_25s_0_pp_2_23, mult_29s_25s_0_pp_3_24, 
        mult_29s_25s_0_pp_3_23, co_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_25, 
        s_mult_29s_25s_0_1_26, mult_29s_25s_0_pp_2_26, mult_29s_25s_0_pp_2_25, 
        mult_29s_25s_0_pp_3_26, mult_29s_25s_0_pp_3_25, s_mult_29s_25s_0_1_27, 
        s_mult_29s_25s_0_1_28, mult_29s_25s_0_pp_2_28, mult_29s_25s_0_pp_2_27, 
        mult_29s_25s_0_pp_3_28, mult_29s_25s_0_pp_3_27, co_mult_29s_25s_0_2_1, 
        s_mult_29s_25s_0_2_10, mult_29s_25s_0_pp_4_10, co_mult_29s_25s_0_2_2, 
        s_mult_29s_25s_0_2_12, s_mult_29s_25s_0_2_11, mult_29s_25s_0_pp_4_12, 
        mult_29s_25s_0_pp_4_11, mult_29s_25s_0_pp_5_12, mult_29s_25s_0_pp_5_11, 
        co_mult_29s_25s_0_2_3, s_mult_29s_25s_0_2_13, s_mult_29s_25s_0_2_14, 
        mult_29s_25s_0_pp_4_14, mult_29s_25s_0_pp_4_13, mult_29s_25s_0_pp_5_14, 
        mult_29s_25s_0_pp_5_13, co_mult_29s_25s_0_2_4, s_mult_29s_25s_0_2_15, 
        s_mult_29s_25s_0_2_16, mult_29s_25s_0_pp_4_16, mult_29s_25s_0_pp_4_15, 
        mult_29s_25s_0_pp_5_16, mult_29s_25s_0_pp_5_15, co_mult_29s_25s_0_2_5, 
        s_mult_29s_25s_0_2_17, s_mult_29s_25s_0_2_18, mult_29s_25s_0_pp_4_18, 
        mult_29s_25s_0_pp_4_17, mult_29s_25s_0_pp_5_18, mult_29s_25s_0_pp_5_17, 
        co_mult_29s_25s_0_2_6, s_mult_29s_25s_0_2_19, s_mult_29s_25s_0_2_20, 
        mult_29s_25s_0_pp_4_20, mult_29s_25s_0_pp_4_19, mult_29s_25s_0_pp_5_20, 
        mult_29s_25s_0_pp_5_19, co_mult_29s_25s_0_2_7, s_mult_29s_25s_0_2_21, 
        s_mult_29s_25s_0_2_22, mult_29s_25s_0_pp_4_22, mult_29s_25s_0_pp_4_21, 
        mult_29s_25s_0_pp_5_22, mult_29s_25s_0_pp_5_21, co_mult_29s_25s_0_2_8, 
        s_mult_29s_25s_0_2_23, s_mult_29s_25s_0_2_24, mult_29s_25s_0_pp_4_24, 
        mult_29s_25s_0_pp_4_23, mult_29s_25s_0_pp_5_24, mult_29s_25s_0_pp_5_23, 
        co_mult_29s_25s_0_2_9, s_mult_29s_25s_0_2_25, s_mult_29s_25s_0_2_26, 
        mult_29s_25s_0_pp_4_26, mult_29s_25s_0_pp_4_25, mult_29s_25s_0_pp_5_26, 
        mult_29s_25s_0_pp_5_25, s_mult_29s_25s_0_2_27, s_mult_29s_25s_0_2_28, 
        mult_29s_25s_0_pp_4_28, mult_29s_25s_0_pp_4_27, mult_29s_25s_0_pp_5_28, 
        mult_29s_25s_0_pp_5_27, co_mult_29s_25s_0_3_1, s_mult_29s_25s_0_3_14, 
        mult_29s_25s_0_pp_6_14, co_mult_29s_25s_0_3_2, s_mult_29s_25s_0_3_15, 
        s_mult_29s_25s_0_3_16, mult_29s_25s_0_pp_6_16, mult_29s_25s_0_pp_6_15, 
        mult_29s_25s_0_pp_7_16, mult_29s_25s_0_pp_7_15, co_mult_29s_25s_0_3_3, 
        s_mult_29s_25s_0_3_17, s_mult_29s_25s_0_3_18, mult_29s_25s_0_pp_6_18, 
        mult_29s_25s_0_pp_6_17, mult_29s_25s_0_pp_7_18, mult_29s_25s_0_pp_7_17, 
        co_mult_29s_25s_0_3_4, s_mult_29s_25s_0_3_19, s_mult_29s_25s_0_3_20, 
        mult_29s_25s_0_pp_6_20, mult_29s_25s_0_pp_6_19, mult_29s_25s_0_pp_7_20, 
        mult_29s_25s_0_pp_7_19, co_mult_29s_25s_0_3_5, s_mult_29s_25s_0_3_21, 
        s_mult_29s_25s_0_3_22, mult_29s_25s_0_pp_6_22, mult_29s_25s_0_pp_6_21, 
        mult_29s_25s_0_pp_7_22, mult_29s_25s_0_pp_7_21, co_mult_29s_25s_0_3_6, 
        s_mult_29s_25s_0_3_23, s_mult_29s_25s_0_3_24, mult_29s_25s_0_pp_6_24, 
        mult_29s_25s_0_pp_6_23, mult_29s_25s_0_pp_7_24, mult_29s_25s_0_pp_7_23, 
        co_mult_29s_25s_0_3_7, s_mult_29s_25s_0_3_25, s_mult_29s_25s_0_3_26, 
        mult_29s_25s_0_pp_6_26, mult_29s_25s_0_pp_6_25, mult_29s_25s_0_pp_7_26, 
        mult_29s_25s_0_pp_7_25, s_mult_29s_25s_0_3_27, s_mult_29s_25s_0_3_28, 
        mult_29s_25s_0_pp_6_28, mult_29s_25s_0_pp_6_27, mult_29s_25s_0_pp_7_28, 
        mult_29s_25s_0_pp_7_27, co_mult_29s_25s_0_4_1, s_mult_29s_25s_0_4_18, 
        mult_29s_25s_0_pp_8_18, co_mult_29s_25s_0_4_2, s_mult_29s_25s_0_4_20, 
        s_mult_29s_25s_0_4_19, mult_29s_25s_0_pp_8_20, mult_29s_25s_0_pp_8_19, 
        mult_29s_25s_0_pp_9_20, mult_29s_25s_0_pp_9_19, co_mult_29s_25s_0_4_3, 
        s_mult_29s_25s_0_4_21, s_mult_29s_25s_0_4_22, mult_29s_25s_0_pp_8_22, 
        mult_29s_25s_0_pp_8_21, mult_29s_25s_0_pp_9_22, mult_29s_25s_0_pp_9_21, 
        co_mult_29s_25s_0_4_4, s_mult_29s_25s_0_4_23, s_mult_29s_25s_0_4_24, 
        mult_29s_25s_0_pp_8_24, mult_29s_25s_0_pp_8_23, mult_29s_25s_0_pp_9_24, 
        mult_29s_25s_0_pp_9_23, co_mult_29s_25s_0_4_5, s_mult_29s_25s_0_4_25, 
        s_mult_29s_25s_0_4_26, mult_29s_25s_0_pp_8_26, mult_29s_25s_0_pp_8_25, 
        mult_29s_25s_0_pp_9_26, mult_29s_25s_0_pp_9_25, s_mult_29s_25s_0_4_27, 
        s_mult_29s_25s_0_4_28, mult_29s_25s_0_pp_8_28, mult_29s_25s_0_pp_8_27, 
        mult_29s_25s_0_pp_9_28, mult_29s_25s_0_pp_9_27, co_mult_29s_25s_0_5_1, 
        s_mult_29s_25s_0_5_22, mult_29s_25s_0_pp_10_22, co_mult_29s_25s_0_5_2, 
        s_mult_29s_25s_0_5_23, s_mult_29s_25s_0_5_24, mult_29s_25s_0_pp_10_24, 
        mult_29s_25s_0_pp_10_23, mult_29s_25s_0_pp_11_24, mult_29s_25s_0_pp_11_23, 
        co_mult_29s_25s_0_5_3, s_mult_29s_25s_0_5_25, s_mult_29s_25s_0_5_26, 
        mult_29s_25s_0_pp_10_26, mult_29s_25s_0_pp_10_25, mult_29s_25s_0_pp_11_26, 
        mult_29s_25s_0_pp_11_25, s_mult_29s_25s_0_5_27, s_mult_29s_25s_0_5_28, 
        mult_29s_25s_0_pp_10_28, mult_29s_25s_0_pp_10_27, mult_29s_25s_0_pp_11_28, 
        mult_29s_25s_0_pp_11_27, co_mult_29s_25s_0_6_1, s_mult_29s_25s_0_6_24, 
        co_mult_29s_25s_0_6_2, s_mult_29s_25s_0_6_25, s_mult_29s_25s_0_6_26, 
        s_mult_29s_25s_0_6_27, s_mult_29s_25s_0_6_28, n21508, n4147, 
        co_mult_29s_25s_0_7_1, co_mult_29s_25s_0_7_2, mult_29s_25s_0_pp_2_5, 
        co_mult_29s_25s_0_7_3, s_mult_29s_25s_0_7_8, co_mult_29s_25s_0_7_4, 
        s_mult_29s_25s_0_7_9, s_mult_29s_25s_0_7_10, co_mult_29s_25s_0_7_5, 
        s_mult_29s_25s_0_7_11, s_mult_29s_25s_0_7_12, co_mult_29s_25s_0_7_6, 
        s_mult_29s_25s_0_7_13, s_mult_29s_25s_0_7_14, co_mult_29s_25s_0_7_7, 
        s_mult_29s_25s_0_7_15, s_mult_29s_25s_0_7_16, co_mult_29s_25s_0_7_8, 
        s_mult_29s_25s_0_7_17, s_mult_29s_25s_0_7_18, co_mult_29s_25s_0_7_9, 
        s_mult_29s_25s_0_7_19, s_mult_29s_25s_0_7_20, co_mult_29s_25s_0_7_10, 
        s_mult_29s_25s_0_7_21, s_mult_29s_25s_0_7_22, co_mult_29s_25s_0_7_11, 
        s_mult_29s_25s_0_7_23, s_mult_29s_25s_0_7_24, co_mult_29s_25s_0_7_12, 
        s_mult_29s_25s_0_7_25, s_mult_29s_25s_0_7_26, s_mult_29s_25s_0_7_27, 
        s_mult_29s_25s_0_7_28, co_mult_29s_25s_0_8_1, s_mult_29s_25s_0_8_12, 
        co_mult_29s_25s_0_8_2, s_mult_29s_25s_0_8_13, s_mult_29s_25s_0_8_14, 
        mult_29s_25s_0_pp_6_13, co_mult_29s_25s_0_8_3, s_mult_29s_25s_0_8_15, 
        s_mult_29s_25s_0_8_16, co_mult_29s_25s_0_8_4, s_mult_29s_25s_0_8_17, 
        s_mult_29s_25s_0_8_18, co_mult_29s_25s_0_8_5, s_mult_29s_25s_0_8_19, 
        s_mult_29s_25s_0_8_20, co_mult_29s_25s_0_8_6, s_mult_29s_25s_0_8_21, 
        s_mult_29s_25s_0_8_22, co_mult_29s_25s_0_8_7, s_mult_29s_25s_0_8_23, 
        s_mult_29s_25s_0_8_24, co_mult_29s_25s_0_8_8, s_mult_29s_25s_0_8_25, 
        s_mult_29s_25s_0_8_26, s_mult_29s_25s_0_8_27, s_mult_29s_25s_0_8_28, 
        co_mult_29s_25s_0_9_1, s_mult_29s_25s_0_9_20, co_mult_29s_25s_0_9_2, 
        s_mult_29s_25s_0_9_21, s_mult_29s_25s_0_9_22, mult_29s_25s_0_pp_10_21, 
        co_mult_29s_25s_0_9_3, s_mult_29s_25s_0_9_24, s_mult_29s_25s_0_9_23, 
        co_mult_29s_25s_0_9_4, s_mult_29s_25s_0_9_25, s_mult_29s_25s_0_9_26, 
        s_mult_29s_25s_0_9_27, s_mult_29s_25s_0_9_28, co_mult_29s_25s_0_10_1, 
        co_mult_29s_25s_0_10_2, mult_29s_25s_0_pp_4_9, co_mult_29s_25s_0_10_3, 
        co_mult_29s_25s_0_10_4, co_mult_29s_25s_0_10_5, s_mult_29s_25s_0_10_16, 
        co_mult_29s_25s_0_10_6, s_mult_29s_25s_0_10_17, s_mult_29s_25s_0_10_18, 
        co_mult_29s_25s_0_10_7, s_mult_29s_25s_0_10_19, s_mult_29s_25s_0_10_20, 
        co_mult_29s_25s_0_10_8, s_mult_29s_25s_0_10_21, s_mult_29s_25s_0_10_22, 
        co_mult_29s_25s_0_10_9, s_mult_29s_25s_0_10_23, s_mult_29s_25s_0_10_24, 
        co_mult_29s_25s_0_10_10, s_mult_29s_25s_0_10_25, s_mult_29s_25s_0_10_26, 
        s_mult_29s_25s_0_10_27, s_mult_29s_25s_0_10_28, co_mult_29s_25s_0_11_1, 
        s_mult_29s_25s_0_11_24, co_mult_29s_25s_0_11_2, s_mult_29s_25s_0_11_25, 
        s_mult_29s_25s_0_11_26, s_mult_29s_25s_0_11_27, s_mult_29s_25s_0_11_28, 
        co_t_mult_29s_25s_0_12_1, co_t_mult_29s_25s_0_12_2, mult_29s_25s_0_pp_8_17, 
        co_t_mult_29s_25s_0_12_3, co_t_mult_29s_25s_0_12_4, co_t_mult_29s_25s_0_12_5, 
        co_t_mult_29s_25s_0_12_6, mult_29s_25s_0_cin_lr_0, mco, mco_1, 
        mco_2, mco_3, mco_4, mco_5, mco_6, mco_7, mco_8, mco_9, 
        mco_10, mco_11, mco_12, mco_14, mco_15, mco_16, mco_17, 
        mco_18, mco_19, mco_20, mco_21, mco_22, mco_23, mco_24, 
        mco_25, mco_28, mco_29, mco_30, mco_31, mco_32, mco_33, 
        mco_34, mco_35, mco_36, mco_37, mco_38, mco_42, mco_43, 
        mco_44, mco_45, mco_46, mco_47, mco_48, mco_49, mco_50, 
        mco_51, mco_56, mco_57, mco_58, mco_59, mco_60, mco_61, 
        mco_62, mco_63, mco_64;
    wire [15:0]n1187;
    
    wire n30, n18815, mco_70, mco_71, mco_72, mco_73, mco_74, 
        mco_75, mco_76, mco_77, mco_84, mco_85, mco_86, mco_87, 
        mco_88, mco_89, mco_90, mco_98, mco_99, mco_100, mco_101, 
        mco_102, mco_103, mco_112, mco_113, mco_114, mco_115, mco_116, 
        mco_126, mco_127, mco_128, mco_129, mco_140, mco_141, mco_142, 
        n21510, n21526, n21543, n20579, mco_154, mco_155, n21520;
    wire [28:0]addIn2_28__N_1337;
    
    wire n5109, n5067, n5157, n5107, n5065, n5155, n5105, n5063, 
        n5153;
    wire [28:0]n121;
    
    wire n5103, n5061, n5151, n5101, n5059, n5149, n5099, n5057, 
        n5147, n5097, n5055, n5145;
    wire [20:0]subIn2_24__N_1301;
    wire [19:0]n3690;
    
    wire n14_adj_1830, n10_adj_1831, n18864, n5095, n5053, n5143, 
        n5093, n5051, n5141, n6_adj_1832, n18865, n5091, n5049, 
        n5139, n5047, n5045, n5137, n19740, n21565, n30_adj_1833;
    wire [15:0]n1166;
    wire [9:0]n2164;
    wire [9:0]n1302;
    
    wire n21528, n15941, n16618;
    wire [9:0]n1346;
    
    wire n9, n7_c;
    wire [15:0]n1208;
    
    wire n30_adj_1834, n10_adj_1835, n8, n4;
    wire [21:0]n2484;
    
    wire n5689, n12666, n5691;
    wire [9:0]n2188;
    wire [9:0]n1390;
    
    wire n21577, n56, n21488, n57, n21583, n21584, n18638;
    wire [24:0]subIn2;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(83[9:15])
    
    wire n16648, n16541, n5701, n5703;
    wire [24:0]n27;
    
    wire n18639, n21569, n18707, n19776, n5693, n19779, n21601, 
        n5695, n19897, n21548, n21552, n18637, n5697, n5699, n18636, 
        n21609, n21529;
    wire [28:0]n588;
    
    wire n21607, n21608, n12641, n5705, n5707, n5709, n5711, n5713, 
        n18706, n5715, n18705, n5717, n5719, n5721, n21509, n21489, 
        n5723, n21490, n21485, n21553;
    wire [20:0]subIn2_24__N_1114;
    
    wire n5725, n18443, n18444, n18635, n5254, n18704, n5729;
    wire [28:0]n618;
    
    wire n20447;
    wire [28:0]addIn2_28__N_1207;
    
    wire n18570, n18442, n18411, n18410, n18409, n18408, n18407, 
        n18406, n18405, n18404, n18400;
    wire [15:0]n1145;
    wire [9:0]n2152;
    
    wire n18401, n18402, n18403, n18399, n18569, n18568, n18703, 
        n18567, n18566, n18702, n18441, n18701, n18700, n18516, 
        n18515, n18514, n18513, n18565, n18440, n18564, n18699, 
        n18563, n18562, n18698, n18512, n18697, n18439, n18561, 
        n18859, n18860, n18696, n18560, n21530, n21491, n18695, 
        n18694, n18559, n18511, n18510, n18558, n18557, n18509, 
        n18438, n18437, n18693, n18692, n18691, n18690, n18508, 
        n21599, n18507, n21487, n18436, n18435, n18689, n12648, 
        n12639, n19668, n18688, n18506, n18434, n18687, n18686, 
        n18685, n18433, n18505, n18684, n18504, n18683, n18432, 
        n18431, n18503, n18502, n18430, n18501, n16636, n18429, 
        n18682, n49, n18681, n18680, n18679, n18428, n18427, n18678, 
        n18677, n18500, n18499, n18498, n18426, n18425, n18497, 
        n18496, n18495, n18424, n18423, n18676, n18675, n18674, 
        n18494, n21610, n18422;
    wire [9:0]n1258;
    
    wire n18421, n18673, n18493, n18492, n18420, n14_adj_1837, n10_adj_1838, 
        n30_adj_1839, n18419, n18491, n18418, n18672, n18671, n18417, 
        n18670, n18416, n18490, n18415, n21486, n19788, n18669, 
        n19732, n18668, n18667, n18666, n18414, n18665, n18664, 
        n18663, n18593, n18592, n18591, n18590, n18589, n18588, 
        n18587, n9_adj_1840, n7_adj_1841, n18586, n18585, n10_adj_1842, 
        n8_adj_1843, n4_adj_1844, n18584, n18645, n18644, n18446, 
        n18445, n18643, n18642, n18641, n18640, n6_adj_1845, n9_adj_1846, 
        n7_adj_1847, n18717, n18716, n10_adj_1848, n18715, n18714, 
        n18713, n8_adj_1849, n4_adj_1850, n9_adj_1851, n7_adj_1852, 
        n10_adj_1853, n8_adj_1854, n4_adj_1855;
    
    FD1P3AX backOut0_i0_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i0.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i0.GSR = "DISABLED";
    FD1S3AX multOut_i0 (.D(multOut_28__N_1178[0]), .CK(clk_N_683), .Q(multOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i0.GSR = "ENABLED";
    FD1P3AX intgOut0_i0 (.D(intgOut1_28__N_766[0]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i0.GSR = "ENABLED";
    FD1P3AX intgOut1_i0 (.D(intgOut1_28__N_766[0]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i0.GSR = "ENABLED";
    FD1P3AX intgOut2_i0 (.D(intgOut1_28__N_766[0]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i0.GSR = "ENABLED";
    FD1P3AX intgOut3_i0 (.D(intgOut1_28__N_766[0]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i0.GSR = "ENABLED";
    FD1P3AX Out0_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i0.GSR = "ENABLED";
    FD1P3AX Out1_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i0.GSR = "ENABLED";
    FD1P3AX Out2_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i0.GSR = "ENABLED";
    FD1P3AX Out3_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i0.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i0.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i0 (.D(backOut1_28__N_1445[0]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i0.GSR = "DISABLED";
    CCU2D add_15798_12 (.A0(addOut[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18711), .COUT(n18712));
    defparam add_15798_12.INIT0 = 16'h5aaa;
    defparam add_15798_12.INIT1 = 16'h5aaa;
    defparam add_15798_12.INJECT1_0 = "NO";
    defparam add_15798_12.INJECT1_1 = "NO";
    FD1S3AX subOut_i0 (.D(subOut_24__N_1135[0]), .CK(clk_N_683), .Q(subOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i0.GSR = "ENABLED";
    CCU2D add_15798_10 (.A0(addOut[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18710), .COUT(n18711));
    defparam add_15798_10.INIT0 = 16'h5555;
    defparam add_15798_10.INIT1 = 16'h5aaa;
    defparam add_15798_10.INJECT1_0 = "NO";
    defparam add_15798_10.INJECT1_1 = "NO";
    FD1P3AX backOut1_i0_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i15.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i0 (.D(n2176[0]), .SP(clk_N_683_enable_392), .CD(n12655), 
            .CK(clk_N_683), .Q(PWMdut_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i0.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i13.GSR = "DISABLED";
    FD1S3IX ss_i2 (.D(n14), .CK(clk_N_683), .CD(ss[4]), .Q(ss[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam ss_i2.GSR = "ENABLED";
    FD1S3IX ss_i3 (.D(n15), .CK(clk_N_683), .CD(ss[4]), .Q(ss[3]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam ss_i3.GSR = "ENABLED";
    FD1S3AY ss_i4 (.D(n19725), .CK(clk_N_683), .Q(ss[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam ss_i4.GSR = "ENABLED";
    FD1P3AX backOut1_i0_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_41), 
            .CK(clk_N_683), .Q(backOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut1_i0_i1.GSR = "DISABLED";
    FD1S3IX ss_i0 (.D(n21572), .CK(clk_N_683), .CD(ss[4]), .Q(ss[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam ss_i0.GSR = "ENABLED";
    FD1S3IX ss_i1 (.D(n21571), .CK(clk_N_683), .CD(ss[4]), .Q(ss[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam ss_i1.GSR = "ENABLED";
    CCU2D add_1179_19 (.A0(n5171), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5173), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18412), 
          .COUT(n18413), .S0(n2244[17]), .S1(n2244[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_19.INIT0 = 16'hf555;
    defparam add_1179_19.INIT1 = 16'hf555;
    defparam add_1179_19.INJECT1_0 = "NO";
    defparam add_1179_19.INJECT1_1 = "NO";
    FD1P3AX dirout_m2_308 (.D(subIn1_24__N_1300), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m2));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dirout_m2_308.GSR = "DISABLED";
    FD1P3AX dirout_m3_309 (.D(dirout_m3_N_1578), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m3));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dirout_m3_309.GSR = "DISABLED";
    FD1P3AX dirout_m1_307 (.D(subIn1_24__N_1113), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m1));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dirout_m1_307.GSR = "DISABLED";
    FD1P3AX dirout_m4_310 (.D(dirout_m4_N_1581), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m4));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dirout_m4_310.GSR = "DISABLED";
    LUT4 i17247_2_lut_3_lut_4_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21554), 
         .D(n21549), .Z(n20450)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam i17247_2_lut_3_lut_4_lut_4_lut.init = 16'hf7e6;
    LUT4 ss_2__bdd_3_lut_rep_313_4_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21550), 
         .D(n21578), .Z(n21522)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(170[9:16])
    defparam ss_2__bdd_3_lut_rep_313_4_lut_4_lut.init = 16'hf7e6;
    LUT4 i1_4_lut_then_4_lut (.A(n22208), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21613)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_else_4_lut (.A(n22208), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21612)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0100;
    LUT4 i17874_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut (.A(n22208), .B(ss[3]), 
         .C(n4138), .D(n21571), .Z(n20179)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17874_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut.init = 16'hf1f0;
    PFUMX mux_1193_i21 (.BLUT(n5129), .ALUT(n5087), .C0(n2436), .Z(n5177));
    LUT4 i3407_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[9]), .C(speed_set_m1[9]), 
         .D(n21500), .Z(n5704)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3407_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n920), .B(n3635), .C(addOut[5]), .D(n22208), 
         .Z(intgOut0_28__N_735[5])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i3393_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[2]), .C(speed_set_m1[2]), 
         .D(n21500), .Z(n5690)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3393_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3395_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[3]), .C(speed_set_m1[3]), 
         .D(n21500), .Z(n5692)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3395_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3397_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[4]), .C(speed_set_m1[4]), 
         .D(n21500), .Z(n5694)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3397_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_139_i1_3_lut (.A(n648[0]), .B(intgOut0[0]), .C(n21551), .Z(n678[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i1_3_lut.init = 16'hcaca;
    LUT4 mux_135_i1_4_lut (.A(backOut2[0]), .B(backOut3[0]), .C(n21524), 
         .D(n15859), .Z(n558[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i1_4_lut.init = 16'hca0a;
    LUT4 mux_139_i5_3_lut (.A(n648[4]), .B(intgOut0[4]), .C(n21551), .Z(n678[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i5_3_lut.init = 16'hcaca;
    LUT4 mux_135_i5_4_lut (.A(backOut2[4]), .B(backOut3[4]), .C(n21524), 
         .D(n15859), .Z(n558[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i5_4_lut.init = 16'hca0a;
    PFUMX mux_1193_i20 (.BLUT(n5127), .ALUT(n5085), .C0(n2436), .Z(n5175));
    LUT4 i3399_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[5]), .C(speed_set_m1[5]), 
         .D(n21500), .Z(n5696)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3399_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3401_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[6]), .C(speed_set_m1[6]), 
         .D(n21500), .Z(n5698)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3401_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3409_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[10]), .C(speed_set_m1[10]), 
         .D(n21500), .Z(n5706)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3409_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3411_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[11]), .C(speed_set_m1[11]), 
         .D(n21500), .Z(n5708)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3411_3_lut_4_lut_4_lut.init = 16'hd8cc;
    PFUMX mux_1193_i19 (.BLUT(n5125), .ALUT(n5083), .C0(n2436), .Z(n5173));
    LUT4 mux_139_i4_3_lut (.A(n648[3]), .B(intgOut0[3]), .C(n21551), .Z(n678[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i4_3_lut.init = 16'hcaca;
    LUT4 mux_135_i4_4_lut (.A(backOut2[3]), .B(backOut3[3]), .C(n21524), 
         .D(n15859), .Z(n558[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i4_4_lut.init = 16'hca0a;
    PFUMX mux_1193_i18 (.BLUT(n5123), .ALUT(n5081), .C0(n2436), .Z(n5171));
    LUT4 i7_4_lut (.A(Out2[3]), .B(n14_adj_1826), .C(n10), .D(Out2[4]), 
         .Z(n18862)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i3413_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[12]), .C(speed_set_m1[12]), 
         .D(n21500), .Z(n5710)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3413_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i6_4_lut (.A(Out2[11]), .B(Out2[7]), .C(Out2[2]), .D(Out2[10]), 
         .Z(n14_adj_1826)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 mux_139_i3_3_lut (.A(n648[2]), .B(intgOut0[2]), .C(n21551), .Z(n678[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i3_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut (.A(Out2[9]), .B(Out2[1]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3415_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[13]), .C(speed_set_m1[13]), 
         .D(n21500), .Z(n5712)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3415_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i4_4_lut (.A(Out2[5]), .B(Out2[6]), .C(Out2[0]), .D(n6), .Z(n18863)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam i4_4_lut.init = 16'hfffe;
    PFUMX mux_1193_i17 (.BLUT(n5121), .ALUT(n5079), .C0(n2436), .Z(n5169));
    LUT4 mux_135_i3_4_lut (.A(backOut2[2]), .B(backOut3[2]), .C(n21524), 
         .D(n15859), .Z(n558[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i3_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut (.A(Out2[8]), .B(Out2[12]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mux_139_i16_3_lut (.A(n648[15]), .B(intgOut0[15]), .C(n21551), 
         .Z(n678[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i16_3_lut.init = 16'hcaca;
    LUT4 mux_135_i16_4_lut (.A(backOut2[15]), .B(backOut3[15]), .C(n21524), 
         .D(n15859), .Z(n558[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i16_4_lut.init = 16'hca0a;
    LUT4 mux_139_i15_3_lut (.A(n648[14]), .B(intgOut0[14]), .C(n21551), 
         .Z(n678[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i15_3_lut.init = 16'hcaca;
    LUT4 i3431_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[20]), .C(speed_set_m1[20]), 
         .D(n21500), .Z(n5728)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3431_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_135_i15_4_lut (.A(backOut2[14]), .B(backOut3[14]), .C(n21524), 
         .D(n15859), .Z(n558[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i15_4_lut.init = 16'hca0a;
    LUT4 i3417_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[14]), .C(speed_set_m1[14]), 
         .D(n21500), .Z(n5714)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3417_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i2959_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[0]), .C(speed_set_m1[0]), 
         .D(n21500), .Z(n5253)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i2959_3_lut_4_lut_4_lut.init = 16'hd8cc;
    PFUMX mux_1193_i16 (.BLUT(n5119), .ALUT(n5077), .C0(n2436), .Z(n5167));
    LUT4 i3391_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[1]), .C(speed_set_m1[1]), 
         .D(n21500), .Z(n5688)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3391_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3423_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[17]), .C(speed_set_m1[17]), 
         .D(n21500), .Z(n5720)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3423_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3405_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[8]), .C(speed_set_m1[8]), 
         .D(n21500), .Z(n5702)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3405_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3403_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[7]), .C(speed_set_m1[7]), 
         .D(n21500), .Z(n5700)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3403_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3419_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[15]), .C(speed_set_m1[15]), 
         .D(n21500), .Z(n5716)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3419_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3421_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[16]), .C(speed_set_m1[16]), 
         .D(n21500), .Z(n5718)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3421_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i3425_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[18]), .C(speed_set_m1[18]), 
         .D(n21500), .Z(n5722)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3425_3_lut_4_lut_4_lut.init = 16'hd8cc;
    PFUMX mux_1193_i15 (.BLUT(n5117), .ALUT(n5075), .C0(n2436), .Z(n5165));
    LUT4 mux_139_i24_3_lut (.A(n648[23]), .B(intgOut0[23]), .C(n21551), 
         .Z(n678[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i24_3_lut.init = 16'hcaca;
    LUT4 n11060_bdd_4_lut (.A(n22196), .B(ss[0]), .C(n22199), .D(ss[1]), 
         .Z(n4138)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam n11060_bdd_4_lut.init = 16'h0410;
    LUT4 mux_135_i24_4_lut (.A(backOut2[23]), .B(backOut3[23]), .C(n21524), 
         .D(n15859), .Z(n558[23])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i24_4_lut.init = 16'hca0a;
    LUT4 i13920_4_lut_4_lut (.A(n920), .B(n3635), .C(addOut[9]), .D(n22208), 
         .Z(intgOut0_28__N_735[9])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13920_4_lut_4_lut.init = 16'h00ba;
    LUT4 i14362_2_lut_rep_275_2_lut_3_lut_4_lut_4_lut (.A(n35), .B(n21500), 
         .C(n42), .D(n21499), .Z(n21484)) /* synthesis lut_function=(A (C+(D))+!A !(B+!(C+(D)))) */ ;
    defparam i14362_2_lut_rep_275_2_lut_3_lut_4_lut_4_lut.init = 16'hbbb0;
    LUT4 mux_139_i23_3_lut (.A(n648[22]), .B(intgOut0[22]), .C(n21551), 
         .Z(n678[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i23_3_lut.init = 16'hcaca;
    LUT4 i3427_3_lut_4_lut_4_lut (.A(n35), .B(speed_set_m2[19]), .C(speed_set_m1[19]), 
         .D(n21500), .Z(n5724)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i3427_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_135_i23_4_lut (.A(backOut2[22]), .B(backOut3[22]), .C(n21524), 
         .D(n15859), .Z(n558[22])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i23_4_lut.init = 16'hca0a;
    CCU2D add_15798_8 (.A0(addOut[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18709), .COUT(n18710));
    defparam add_15798_8.INIT0 = 16'h5555;
    defparam add_15798_8.INIT1 = 16'h5aaa;
    defparam add_15798_8.INJECT1_0 = "NO";
    defparam add_15798_8.INJECT1_1 = "NO";
    LUT4 i14363_1_lut_rep_274_2_lut_2_lut_3_lut_4_lut_4_lut (.A(n35), .B(n21500), 
         .C(n42), .D(n21499), .Z(n21483)) /* synthesis lut_function=(!(A (C+(D))+!A !(B+!(C+(D))))) */ ;
    defparam i14363_1_lut_rep_274_2_lut_2_lut_3_lut_4_lut_4_lut.init = 16'h444f;
    PFUMX mux_1193_i14 (.BLUT(n5115), .ALUT(n5073), .C0(n2436), .Z(n5163));
    LUT4 mux_139_i2_3_lut (.A(n648[1]), .B(intgOut0[1]), .C(n21551), .Z(n678[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_43 (.A(n920), .B(n3635), .C(addOut[1]), 
         .D(n22208), .Z(intgOut0_28__N_735[1])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_43.init = 16'h0010;
    LUT4 mux_135_i2_4_lut (.A(backOut2[1]), .B(backOut3[1]), .C(n21524), 
         .D(n15859), .Z(n558[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i2_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_3_lut_4_lut_adj_44 (.A(n920), .B(n3635), .C(addOut[0]), 
         .D(n22208), .Z(intgOut1_28__N_766[0])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_44.init = 16'h0010;
    PFUMX mux_1193_i13 (.BLUT(n5113), .ALUT(n5071), .C0(n2436), .Z(n5161));
    CCU2D add_15798_6 (.A0(addOut[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18708), .COUT(n18709));
    defparam add_15798_6.INIT0 = 16'h5555;
    defparam add_15798_6.INIT1 = 16'h5555;
    defparam add_15798_6.INJECT1_0 = "NO";
    defparam add_15798_6.INJECT1_1 = "NO";
    LUT4 mux_139_i14_3_lut (.A(n648[13]), .B(intgOut0[13]), .C(n21551), 
         .Z(n678[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i14_3_lut.init = 16'hcaca;
    LUT4 mux_135_i14_4_lut (.A(backOut2[13]), .B(backOut3[13]), .C(n21524), 
         .D(n15859), .Z(n558[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i14_4_lut.init = 16'hca0a;
    LUT4 mux_139_i13_3_lut (.A(n648[12]), .B(intgOut0[12]), .C(n21551), 
         .Z(n678[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i13_3_lut.init = 16'hcaca;
    LUT4 mux_135_i13_4_lut (.A(backOut2[12]), .B(backOut3[12]), .C(n21524), 
         .D(n15859), .Z(n558[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i13_4_lut.init = 16'hca0a;
    LUT4 i7_4_lut_adj_45 (.A(Out1[3]), .B(n14_adj_1827), .C(n10_adj_1828), 
         .D(Out1[4]), .Z(n18821)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam i7_4_lut_adj_45.init = 16'hfffe;
    LUT4 i6_4_lut_adj_46 (.A(Out1[11]), .B(Out1[7]), .C(Out1[2]), .D(Out1[10]), 
         .Z(n14_adj_1827)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam i6_4_lut_adj_46.init = 16'hfffe;
    LUT4 i2_2_lut_adj_47 (.A(Out1[9]), .B(Out1[1]), .Z(n10_adj_1828)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam i2_2_lut_adj_47.init = 16'heeee;
    LUT4 mux_139_i22_3_lut (.A(n648[21]), .B(intgOut0[21]), .C(n21551), 
         .Z(n678[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i22_3_lut.init = 16'hcaca;
    PFUMX mux_1193_i12 (.BLUT(n5111), .ALUT(n5069), .C0(n2436), .Z(n5159));
    LUT4 mux_135_i22_4_lut (.A(backOut2[21]), .B(backOut3[21]), .C(n21524), 
         .D(n15859), .Z(n558[21])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i22_4_lut.init = 16'hca0a;
    LUT4 i4_4_lut_adj_48 (.A(Out1[5]), .B(Out1[6]), .C(Out1[0]), .D(n6_adj_1829), 
         .Z(n18822)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam i4_4_lut_adj_48.init = 16'hfffe;
    LUT4 mux_139_i12_3_lut (.A(n648[11]), .B(intgOut0[11]), .C(n21551), 
         .Z(n678[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i12_3_lut.init = 16'hcaca;
    LUT4 mux_135_i12_4_lut (.A(backOut2[11]), .B(backOut3[11]), .C(n21524), 
         .D(n15859), .Z(n558[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i12_4_lut.init = 16'hca0a;
    LUT4 mux_139_i21_3_lut (.A(n648[20]), .B(intgOut0[20]), .C(n21551), 
         .Z(n678[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i21_3_lut.init = 16'hcaca;
    AND2 AND2_t64 (.A(subOut[0]), .B(GND_net), .Z(multOut_28__N_1178[0])) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1256[10:66])
    AND2 AND2_t61 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1262[10:66])
    AND2 AND2_t58 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1268[10:66])
    AND2 AND2_t55 (.A(subOut[0]), .B(multIn2[6]), .Z(mult_29s_25s_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1274[10:66])
    LUT4 mux_135_i21_4_lut (.A(backOut2[20]), .B(backOut3[20]), .C(n21524), 
         .D(n15859), .Z(n558[20])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i21_4_lut.init = 16'hca0a;
    AND2 AND2_t52 (.A(subOut[0]), .B(multIn2[6]), .Z(mult_29s_25s_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1280[10:66])
    LUT4 mux_139_i29_3_lut (.A(n648[28]), .B(intgOut0[28]), .C(n21551), 
         .Z(n678[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i29_3_lut.init = 16'hcaca;
    AND2 AND2_t49 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_5_10)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1286[10:68])
    AND2 AND2_t46 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_6_12)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1292[10:68])
    AND2 AND2_t43 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_7_14)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1298[10:68])
    LUT4 mux_135_i29_4_lut (.A(backOut2[28]), .B(backOut3[28]), .C(n21524), 
         .D(n15859), .Z(n558[28])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i29_4_lut.init = 16'hca0a;
    AND2 AND2_t40 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_8_16)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1304[10:68])
    AND2 AND2_t37 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_9_18)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1310[10:68])
    AND2 AND2_t34 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_10_20)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1316[10:69])
    AND2 AND2_t31 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_11_22)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1322[10:69])
    ND2 ND2_t28 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    ND2 ND2_t27 (.A(subOut[1]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_25)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    ND2 ND2_t26 (.A(subOut[2]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    ND2 ND2_t25 (.A(subOut[3]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_27)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    ND2 ND2_t24 (.A(subOut[4]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 i1_2_lut_adj_49 (.A(Out1[8]), .B(Out1[12]), .Z(n6_adj_1829)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam i1_2_lut_adj_49.init = 16'heeee;
    LUT4 mux_139_i11_3_lut (.A(n648[10]), .B(intgOut0[10]), .C(n21551), 
         .Z(n678[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i11_3_lut.init = 16'hcaca;
    LUT4 i13917_3_lut_4_lut (.A(n920), .B(n3635), .C(n22208), .D(addOut[6]), 
         .Z(intgOut0_28__N_735[6])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i13917_3_lut_4_lut.init = 16'h0f0e;
    LUT4 mux_135_i11_4_lut (.A(backOut2[10]), .B(backOut3[10]), .C(n21524), 
         .D(n15859), .Z(n558[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i11_4_lut.init = 16'hca0a;
    FADD2B mult_29s_25s_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_12 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_14 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_16 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_18 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_20 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_22 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_0_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_0_2), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_1_2), .CI(GND_net), .COUT(co_mult_29s_25s_0_0_1), 
           .S1(multOut_28__N_1178[2])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_2 (.A0(mult_29s_25s_0_pp_0_3), .A1(mult_29s_25s_0_pp_0_4), 
           .B0(mult_29s_25s_0_pp_1_3), .B1(mult_29s_25s_0_pp_1_4), .CI(co_mult_29s_25s_0_0_1), 
           .COUT(co_mult_29s_25s_0_0_2), .S0(multOut_28__N_1178[3]), .S1(s_mult_29s_25s_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_3 (.A0(mult_29s_25s_0_pp_0_5), .A1(mult_29s_25s_0_pp_0_6), 
           .B0(mult_29s_25s_0_pp_1_5), .B1(mult_29s_25s_0_pp_1_6), .CI(co_mult_29s_25s_0_0_2), 
           .COUT(co_mult_29s_25s_0_0_3), .S0(s_mult_29s_25s_0_0_5), .S1(s_mult_29s_25s_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_4 (.A0(mult_29s_25s_0_pp_0_7), .A1(mult_29s_25s_0_pp_0_8), 
           .B0(mult_29s_25s_0_pp_1_7), .B1(mult_29s_25s_0_pp_1_8), .CI(co_mult_29s_25s_0_0_3), 
           .COUT(co_mult_29s_25s_0_0_4), .S0(s_mult_29s_25s_0_0_7), .S1(s_mult_29s_25s_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_5 (.A0(mult_29s_25s_0_pp_0_9), .A1(mult_29s_25s_0_pp_0_10), 
           .B0(mult_29s_25s_0_pp_1_9), .B1(mult_29s_25s_0_pp_1_10), .CI(co_mult_29s_25s_0_0_4), 
           .COUT(co_mult_29s_25s_0_0_5), .S0(s_mult_29s_25s_0_0_9), .S1(s_mult_29s_25s_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_6 (.A0(mult_29s_25s_0_pp_0_11), .A1(mult_29s_25s_0_pp_0_12), 
           .B0(mult_29s_25s_0_pp_1_11), .B1(mult_29s_25s_0_pp_1_12), .CI(co_mult_29s_25s_0_0_5), 
           .COUT(co_mult_29s_25s_0_0_6), .S0(s_mult_29s_25s_0_0_11), .S1(s_mult_29s_25s_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_7 (.A0(mult_29s_25s_0_pp_0_13), .A1(mult_29s_25s_0_pp_0_14), 
           .B0(mult_29s_25s_0_pp_1_13), .B1(mult_29s_25s_0_pp_1_14), .CI(co_mult_29s_25s_0_0_6), 
           .COUT(co_mult_29s_25s_0_0_7), .S0(s_mult_29s_25s_0_0_13), .S1(s_mult_29s_25s_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_8 (.A0(mult_29s_25s_0_pp_0_15), .A1(mult_29s_25s_0_pp_0_16), 
           .B0(mult_29s_25s_0_pp_1_15), .B1(mult_29s_25s_0_pp_1_16), .CI(co_mult_29s_25s_0_0_7), 
           .COUT(co_mult_29s_25s_0_0_8), .S0(s_mult_29s_25s_0_0_15), .S1(s_mult_29s_25s_0_0_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_9 (.A0(mult_29s_25s_0_pp_0_17), .A1(mult_29s_25s_0_pp_0_18), 
           .B0(mult_29s_25s_0_pp_1_17), .B1(mult_29s_25s_0_pp_1_18), .CI(co_mult_29s_25s_0_0_8), 
           .COUT(co_mult_29s_25s_0_0_9), .S0(s_mult_29s_25s_0_0_17), .S1(s_mult_29s_25s_0_0_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_10 (.A0(mult_29s_25s_0_pp_0_19), .A1(mult_29s_25s_0_pp_0_20), 
           .B0(mult_29s_25s_0_pp_1_19), .B1(mult_29s_25s_0_pp_1_20), .CI(co_mult_29s_25s_0_0_9), 
           .COUT(co_mult_29s_25s_0_0_10), .S0(s_mult_29s_25s_0_0_19), .S1(s_mult_29s_25s_0_0_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_11 (.A0(mult_29s_25s_0_pp_0_21), .A1(mult_29s_25s_0_pp_0_22), 
           .B0(mult_29s_25s_0_pp_1_21), .B1(mult_29s_25s_0_pp_1_22), .CI(co_mult_29s_25s_0_0_10), 
           .COUT(co_mult_29s_25s_0_0_11), .S0(s_mult_29s_25s_0_0_21), .S1(s_mult_29s_25s_0_0_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_12 (.A0(mult_29s_25s_0_pp_0_23), .A1(mult_29s_25s_0_pp_0_24), 
           .B0(mult_29s_25s_0_pp_1_23), .B1(mult_29s_25s_0_pp_1_24), .CI(co_mult_29s_25s_0_0_11), 
           .COUT(co_mult_29s_25s_0_0_12), .S0(s_mult_29s_25s_0_0_23), .S1(s_mult_29s_25s_0_0_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_13 (.A0(mult_29s_25s_0_pp_0_25), .A1(mult_29s_25s_0_pp_0_26), 
           .B0(mult_29s_25s_0_pp_1_25), .B1(mult_29s_25s_0_pp_1_26), .CI(co_mult_29s_25s_0_0_12), 
           .COUT(co_mult_29s_25s_0_0_13), .S0(s_mult_29s_25s_0_0_25), .S1(s_mult_29s_25s_0_0_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_14 (.A0(mult_29s_25s_0_pp_0_27), .A1(mult_29s_25s_0_pp_0_28), 
           .B0(mult_29s_25s_0_pp_1_27), .B1(mult_29s_25s_0_pp_1_28), .CI(co_mult_29s_25s_0_0_13), 
           .S0(s_mult_29s_25s_0_0_27), .S1(s_mult_29s_25s_0_0_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_1_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_2_6), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_3_6), .CI(GND_net), .COUT(co_mult_29s_25s_0_1_1), 
           .S1(s_mult_29s_25s_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_2 (.A0(mult_29s_25s_0_pp_2_7), .A1(mult_29s_25s_0_pp_2_8), 
           .B0(mult_29s_25s_0_pp_3_7), .B1(mult_29s_25s_0_pp_3_8), .CI(co_mult_29s_25s_0_1_1), 
           .COUT(co_mult_29s_25s_0_1_2), .S0(s_mult_29s_25s_0_1_7), .S1(s_mult_29s_25s_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_3 (.A0(mult_29s_25s_0_pp_2_9), .A1(mult_29s_25s_0_pp_2_10), 
           .B0(mult_29s_25s_0_pp_3_9), .B1(mult_29s_25s_0_pp_3_10), .CI(co_mult_29s_25s_0_1_2), 
           .COUT(co_mult_29s_25s_0_1_3), .S0(s_mult_29s_25s_0_1_9), .S1(s_mult_29s_25s_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_4 (.A0(mult_29s_25s_0_pp_2_11), .A1(mult_29s_25s_0_pp_2_12), 
           .B0(mult_29s_25s_0_pp_3_11), .B1(mult_29s_25s_0_pp_3_12), .CI(co_mult_29s_25s_0_1_3), 
           .COUT(co_mult_29s_25s_0_1_4), .S0(s_mult_29s_25s_0_1_11), .S1(s_mult_29s_25s_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_5 (.A0(mult_29s_25s_0_pp_2_13), .A1(mult_29s_25s_0_pp_2_14), 
           .B0(mult_29s_25s_0_pp_3_13), .B1(mult_29s_25s_0_pp_3_14), .CI(co_mult_29s_25s_0_1_4), 
           .COUT(co_mult_29s_25s_0_1_5), .S0(s_mult_29s_25s_0_1_13), .S1(s_mult_29s_25s_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_6 (.A0(mult_29s_25s_0_pp_2_15), .A1(mult_29s_25s_0_pp_2_16), 
           .B0(mult_29s_25s_0_pp_3_15), .B1(mult_29s_25s_0_pp_3_16), .CI(co_mult_29s_25s_0_1_5), 
           .COUT(co_mult_29s_25s_0_1_6), .S0(s_mult_29s_25s_0_1_15), .S1(s_mult_29s_25s_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_7 (.A0(mult_29s_25s_0_pp_2_17), .A1(mult_29s_25s_0_pp_2_18), 
           .B0(mult_29s_25s_0_pp_3_17), .B1(mult_29s_25s_0_pp_3_18), .CI(co_mult_29s_25s_0_1_6), 
           .COUT(co_mult_29s_25s_0_1_7), .S0(s_mult_29s_25s_0_1_17), .S1(s_mult_29s_25s_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_8 (.A0(mult_29s_25s_0_pp_2_19), .A1(mult_29s_25s_0_pp_2_20), 
           .B0(mult_29s_25s_0_pp_3_19), .B1(mult_29s_25s_0_pp_3_20), .CI(co_mult_29s_25s_0_1_7), 
           .COUT(co_mult_29s_25s_0_1_8), .S0(s_mult_29s_25s_0_1_19), .S1(s_mult_29s_25s_0_1_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_9 (.A0(mult_29s_25s_0_pp_2_21), .A1(mult_29s_25s_0_pp_2_22), 
           .B0(mult_29s_25s_0_pp_3_21), .B1(mult_29s_25s_0_pp_3_22), .CI(co_mult_29s_25s_0_1_8), 
           .COUT(co_mult_29s_25s_0_1_9), .S0(s_mult_29s_25s_0_1_21), .S1(s_mult_29s_25s_0_1_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_10 (.A0(mult_29s_25s_0_pp_2_23), .A1(mult_29s_25s_0_pp_2_24), 
           .B0(mult_29s_25s_0_pp_3_23), .B1(mult_29s_25s_0_pp_3_24), .CI(co_mult_29s_25s_0_1_9), 
           .COUT(co_mult_29s_25s_0_1_10), .S0(s_mult_29s_25s_0_1_23), .S1(s_mult_29s_25s_0_1_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_11 (.A0(mult_29s_25s_0_pp_2_25), .A1(mult_29s_25s_0_pp_2_26), 
           .B0(mult_29s_25s_0_pp_3_25), .B1(mult_29s_25s_0_pp_3_26), .CI(co_mult_29s_25s_0_1_10), 
           .COUT(co_mult_29s_25s_0_1_11), .S0(s_mult_29s_25s_0_1_25), .S1(s_mult_29s_25s_0_1_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_12 (.A0(mult_29s_25s_0_pp_2_27), .A1(mult_29s_25s_0_pp_2_28), 
           .B0(mult_29s_25s_0_pp_3_27), .B1(mult_29s_25s_0_pp_3_28), .CI(co_mult_29s_25s_0_1_11), 
           .S0(s_mult_29s_25s_0_1_27), .S1(s_mult_29s_25s_0_1_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_139_i10_3_lut (.A(n648[9]), .B(intgOut0[9]), .C(n21551), 
         .Z(n678[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i10_3_lut.init = 16'hcaca;
    FADD2B Cadd_mult_29s_25s_0_2_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_4_10), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_5_10), .CI(GND_net), .COUT(co_mult_29s_25s_0_2_1), 
           .S1(s_mult_29s_25s_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_2 (.A0(mult_29s_25s_0_pp_4_11), .A1(mult_29s_25s_0_pp_4_12), 
           .B0(mult_29s_25s_0_pp_5_11), .B1(mult_29s_25s_0_pp_5_12), .CI(co_mult_29s_25s_0_2_1), 
           .COUT(co_mult_29s_25s_0_2_2), .S0(s_mult_29s_25s_0_2_11), .S1(s_mult_29s_25s_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_3 (.A0(mult_29s_25s_0_pp_4_13), .A1(mult_29s_25s_0_pp_4_14), 
           .B0(mult_29s_25s_0_pp_5_13), .B1(mult_29s_25s_0_pp_5_14), .CI(co_mult_29s_25s_0_2_2), 
           .COUT(co_mult_29s_25s_0_2_3), .S0(s_mult_29s_25s_0_2_13), .S1(s_mult_29s_25s_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_4 (.A0(mult_29s_25s_0_pp_4_15), .A1(mult_29s_25s_0_pp_4_16), 
           .B0(mult_29s_25s_0_pp_5_15), .B1(mult_29s_25s_0_pp_5_16), .CI(co_mult_29s_25s_0_2_3), 
           .COUT(co_mult_29s_25s_0_2_4), .S0(s_mult_29s_25s_0_2_15), .S1(s_mult_29s_25s_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_5 (.A0(mult_29s_25s_0_pp_4_17), .A1(mult_29s_25s_0_pp_4_18), 
           .B0(mult_29s_25s_0_pp_5_17), .B1(mult_29s_25s_0_pp_5_18), .CI(co_mult_29s_25s_0_2_4), 
           .COUT(co_mult_29s_25s_0_2_5), .S0(s_mult_29s_25s_0_2_17), .S1(s_mult_29s_25s_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_6 (.A0(mult_29s_25s_0_pp_4_19), .A1(mult_29s_25s_0_pp_4_20), 
           .B0(mult_29s_25s_0_pp_5_19), .B1(mult_29s_25s_0_pp_5_20), .CI(co_mult_29s_25s_0_2_5), 
           .COUT(co_mult_29s_25s_0_2_6), .S0(s_mult_29s_25s_0_2_19), .S1(s_mult_29s_25s_0_2_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_7 (.A0(mult_29s_25s_0_pp_4_21), .A1(mult_29s_25s_0_pp_4_22), 
           .B0(mult_29s_25s_0_pp_5_21), .B1(mult_29s_25s_0_pp_5_22), .CI(co_mult_29s_25s_0_2_6), 
           .COUT(co_mult_29s_25s_0_2_7), .S0(s_mult_29s_25s_0_2_21), .S1(s_mult_29s_25s_0_2_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_8 (.A0(mult_29s_25s_0_pp_4_23), .A1(mult_29s_25s_0_pp_4_24), 
           .B0(mult_29s_25s_0_pp_5_23), .B1(mult_29s_25s_0_pp_5_24), .CI(co_mult_29s_25s_0_2_7), 
           .COUT(co_mult_29s_25s_0_2_8), .S0(s_mult_29s_25s_0_2_23), .S1(s_mult_29s_25s_0_2_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_9 (.A0(mult_29s_25s_0_pp_4_25), .A1(mult_29s_25s_0_pp_4_26), 
           .B0(mult_29s_25s_0_pp_5_25), .B1(mult_29s_25s_0_pp_5_26), .CI(co_mult_29s_25s_0_2_8), 
           .COUT(co_mult_29s_25s_0_2_9), .S0(s_mult_29s_25s_0_2_25), .S1(s_mult_29s_25s_0_2_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_10 (.A0(mult_29s_25s_0_pp_4_27), .A1(mult_29s_25s_0_pp_4_28), 
           .B0(mult_29s_25s_0_pp_5_27), .B1(mult_29s_25s_0_pp_5_28), .CI(co_mult_29s_25s_0_2_9), 
           .S0(s_mult_29s_25s_0_2_27), .S1(s_mult_29s_25s_0_2_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_135_i10_4_lut (.A(backOut2[9]), .B(backOut3[9]), .C(n21524), 
         .D(n15859), .Z(n558[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i10_4_lut.init = 16'hca0a;
    FADD2B Cadd_mult_29s_25s_0_3_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_6_14), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_7_14), .CI(GND_net), .COUT(co_mult_29s_25s_0_3_1), 
           .S1(s_mult_29s_25s_0_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_2 (.A0(mult_29s_25s_0_pp_6_15), .A1(mult_29s_25s_0_pp_6_16), 
           .B0(mult_29s_25s_0_pp_7_15), .B1(mult_29s_25s_0_pp_7_16), .CI(co_mult_29s_25s_0_3_1), 
           .COUT(co_mult_29s_25s_0_3_2), .S0(s_mult_29s_25s_0_3_15), .S1(s_mult_29s_25s_0_3_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_3 (.A0(mult_29s_25s_0_pp_6_17), .A1(mult_29s_25s_0_pp_6_18), 
           .B0(mult_29s_25s_0_pp_7_17), .B1(mult_29s_25s_0_pp_7_18), .CI(co_mult_29s_25s_0_3_2), 
           .COUT(co_mult_29s_25s_0_3_3), .S0(s_mult_29s_25s_0_3_17), .S1(s_mult_29s_25s_0_3_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_4 (.A0(mult_29s_25s_0_pp_6_19), .A1(mult_29s_25s_0_pp_6_20), 
           .B0(mult_29s_25s_0_pp_7_19), .B1(mult_29s_25s_0_pp_7_20), .CI(co_mult_29s_25s_0_3_3), 
           .COUT(co_mult_29s_25s_0_3_4), .S0(s_mult_29s_25s_0_3_19), .S1(s_mult_29s_25s_0_3_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_5 (.A0(mult_29s_25s_0_pp_6_21), .A1(mult_29s_25s_0_pp_6_22), 
           .B0(mult_29s_25s_0_pp_7_21), .B1(mult_29s_25s_0_pp_7_22), .CI(co_mult_29s_25s_0_3_4), 
           .COUT(co_mult_29s_25s_0_3_5), .S0(s_mult_29s_25s_0_3_21), .S1(s_mult_29s_25s_0_3_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_6 (.A0(mult_29s_25s_0_pp_6_23), .A1(mult_29s_25s_0_pp_6_24), 
           .B0(mult_29s_25s_0_pp_7_23), .B1(mult_29s_25s_0_pp_7_24), .CI(co_mult_29s_25s_0_3_5), 
           .COUT(co_mult_29s_25s_0_3_6), .S0(s_mult_29s_25s_0_3_23), .S1(s_mult_29s_25s_0_3_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_7 (.A0(mult_29s_25s_0_pp_6_25), .A1(mult_29s_25s_0_pp_6_26), 
           .B0(mult_29s_25s_0_pp_7_25), .B1(mult_29s_25s_0_pp_7_26), .CI(co_mult_29s_25s_0_3_6), 
           .COUT(co_mult_29s_25s_0_3_7), .S0(s_mult_29s_25s_0_3_25), .S1(s_mult_29s_25s_0_3_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_8 (.A0(mult_29s_25s_0_pp_6_27), .A1(mult_29s_25s_0_pp_6_28), 
           .B0(mult_29s_25s_0_pp_7_27), .B1(mult_29s_25s_0_pp_7_28), .CI(co_mult_29s_25s_0_3_7), 
           .S0(s_mult_29s_25s_0_3_27), .S1(s_mult_29s_25s_0_3_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_139_i20_3_lut (.A(n648[19]), .B(intgOut0[19]), .C(n21551), 
         .Z(n678[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i20_3_lut.init = 16'hcaca;
    LUT4 mux_135_i20_4_lut (.A(backOut2[19]), .B(backOut3[19]), .C(n21524), 
         .D(n15859), .Z(n558[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i20_4_lut.init = 16'hca0a;
    FADD2B Cadd_mult_29s_25s_0_4_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_8_18), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_9_18), .CI(GND_net), .COUT(co_mult_29s_25s_0_4_1), 
           .S1(s_mult_29s_25s_0_4_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_2 (.A0(mult_29s_25s_0_pp_8_19), .A1(mult_29s_25s_0_pp_8_20), 
           .B0(mult_29s_25s_0_pp_9_19), .B1(mult_29s_25s_0_pp_9_20), .CI(co_mult_29s_25s_0_4_1), 
           .COUT(co_mult_29s_25s_0_4_2), .S0(s_mult_29s_25s_0_4_19), .S1(s_mult_29s_25s_0_4_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_3 (.A0(mult_29s_25s_0_pp_8_21), .A1(mult_29s_25s_0_pp_8_22), 
           .B0(mult_29s_25s_0_pp_9_21), .B1(mult_29s_25s_0_pp_9_22), .CI(co_mult_29s_25s_0_4_2), 
           .COUT(co_mult_29s_25s_0_4_3), .S0(s_mult_29s_25s_0_4_21), .S1(s_mult_29s_25s_0_4_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_4 (.A0(mult_29s_25s_0_pp_8_23), .A1(mult_29s_25s_0_pp_8_24), 
           .B0(mult_29s_25s_0_pp_9_23), .B1(mult_29s_25s_0_pp_9_24), .CI(co_mult_29s_25s_0_4_3), 
           .COUT(co_mult_29s_25s_0_4_4), .S0(s_mult_29s_25s_0_4_23), .S1(s_mult_29s_25s_0_4_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_5 (.A0(mult_29s_25s_0_pp_8_25), .A1(mult_29s_25s_0_pp_8_26), 
           .B0(mult_29s_25s_0_pp_9_25), .B1(mult_29s_25s_0_pp_9_26), .CI(co_mult_29s_25s_0_4_4), 
           .COUT(co_mult_29s_25s_0_4_5), .S0(s_mult_29s_25s_0_4_25), .S1(s_mult_29s_25s_0_4_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_6 (.A0(mult_29s_25s_0_pp_8_27), .A1(mult_29s_25s_0_pp_8_28), 
           .B0(mult_29s_25s_0_pp_9_27), .B1(mult_29s_25s_0_pp_9_28), .CI(co_mult_29s_25s_0_4_5), 
           .S0(s_mult_29s_25s_0_4_27), .S1(s_mult_29s_25s_0_4_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_5_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_10_22), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_11_22), .CI(GND_net), .COUT(co_mult_29s_25s_0_5_1), 
           .S1(s_mult_29s_25s_0_5_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_2 (.A0(mult_29s_25s_0_pp_10_23), .A1(mult_29s_25s_0_pp_10_24), 
           .B0(mult_29s_25s_0_pp_11_23), .B1(mult_29s_25s_0_pp_11_24), .CI(co_mult_29s_25s_0_5_1), 
           .COUT(co_mult_29s_25s_0_5_2), .S0(s_mult_29s_25s_0_5_23), .S1(s_mult_29s_25s_0_5_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_3 (.A0(mult_29s_25s_0_pp_10_25), .A1(mult_29s_25s_0_pp_10_26), 
           .B0(mult_29s_25s_0_pp_11_25), .B1(mult_29s_25s_0_pp_11_26), .CI(co_mult_29s_25s_0_5_2), 
           .COUT(co_mult_29s_25s_0_5_3), .S0(s_mult_29s_25s_0_5_25), .S1(s_mult_29s_25s_0_5_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_4 (.A0(mult_29s_25s_0_pp_10_27), .A1(mult_29s_25s_0_pp_10_28), 
           .B0(mult_29s_25s_0_pp_11_27), .B1(mult_29s_25s_0_pp_11_28), .CI(co_mult_29s_25s_0_5_3), 
           .S0(s_mult_29s_25s_0_5_27), .S1(s_mult_29s_25s_0_5_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_6_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_12_24), 
           .B0(GND_net), .B1(VCC_net), .CI(GND_net), .COUT(co_mult_29s_25s_0_6_1), 
           .S1(s_mult_29s_25s_0_6_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_2 (.A0(mult_29s_25s_0_pp_12_25), .A1(mult_29s_25s_0_pp_12_26), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_1), .COUT(co_mult_29s_25s_0_6_2), 
           .S0(s_mult_29s_25s_0_6_25), .S1(s_mult_29s_25s_0_6_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_3 (.A0(mult_29s_25s_0_pp_12_27), .A1(mult_29s_25s_0_pp_12_28), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_2), .S0(s_mult_29s_25s_0_6_27), 
           .S1(s_mult_29s_25s_0_6_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 i13649_3_lut_4_lut (.A(n21524), .B(n21508), .C(multIn2[6]), .D(n4147), 
         .Z(multIn2[3])) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i13649_3_lut_4_lut.init = 16'hff07;
    LUT4 i13648_3_lut_4_lut (.A(n21524), .B(n21508), .C(multIn2[6]), .D(n4147), 
         .Z(multIn2[5])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;
    defparam i13648_3_lut_4_lut.init = 16'h00f7;
    FADD2B Cadd_mult_29s_25s_0_7_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_0_4), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_2_4), .CI(GND_net), .COUT(co_mult_29s_25s_0_7_1), 
           .S1(multOut_28__N_1178[4])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_2 (.A0(s_mult_29s_25s_0_0_5), .A1(s_mult_29s_25s_0_0_6), 
           .B0(mult_29s_25s_0_pp_2_5), .B1(s_mult_29s_25s_0_1_6), .CI(co_mult_29s_25s_0_7_1), 
           .COUT(co_mult_29s_25s_0_7_2), .S0(multOut_28__N_1178[5]), .S1(multOut_28__N_1178[6])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_3 (.A0(s_mult_29s_25s_0_0_7), .A1(s_mult_29s_25s_0_0_8), 
           .B0(s_mult_29s_25s_0_1_7), .B1(s_mult_29s_25s_0_1_8), .CI(co_mult_29s_25s_0_7_2), 
           .COUT(co_mult_29s_25s_0_7_3), .S0(multOut_28__N_1178[7]), .S1(s_mult_29s_25s_0_7_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_4 (.A0(s_mult_29s_25s_0_0_9), .A1(s_mult_29s_25s_0_0_10), 
           .B0(s_mult_29s_25s_0_1_9), .B1(s_mult_29s_25s_0_1_10), .CI(co_mult_29s_25s_0_7_3), 
           .COUT(co_mult_29s_25s_0_7_4), .S0(s_mult_29s_25s_0_7_9), .S1(s_mult_29s_25s_0_7_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_5 (.A0(s_mult_29s_25s_0_0_11), .A1(s_mult_29s_25s_0_0_12), 
           .B0(s_mult_29s_25s_0_1_11), .B1(s_mult_29s_25s_0_1_12), .CI(co_mult_29s_25s_0_7_4), 
           .COUT(co_mult_29s_25s_0_7_5), .S0(s_mult_29s_25s_0_7_11), .S1(s_mult_29s_25s_0_7_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_6 (.A0(s_mult_29s_25s_0_0_13), .A1(s_mult_29s_25s_0_0_14), 
           .B0(s_mult_29s_25s_0_1_13), .B1(s_mult_29s_25s_0_1_14), .CI(co_mult_29s_25s_0_7_5), 
           .COUT(co_mult_29s_25s_0_7_6), .S0(s_mult_29s_25s_0_7_13), .S1(s_mult_29s_25s_0_7_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_7 (.A0(s_mult_29s_25s_0_0_15), .A1(s_mult_29s_25s_0_0_16), 
           .B0(s_mult_29s_25s_0_1_15), .B1(s_mult_29s_25s_0_1_16), .CI(co_mult_29s_25s_0_7_6), 
           .COUT(co_mult_29s_25s_0_7_7), .S0(s_mult_29s_25s_0_7_15), .S1(s_mult_29s_25s_0_7_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_8 (.A0(s_mult_29s_25s_0_0_17), .A1(s_mult_29s_25s_0_0_18), 
           .B0(s_mult_29s_25s_0_1_17), .B1(s_mult_29s_25s_0_1_18), .CI(co_mult_29s_25s_0_7_7), 
           .COUT(co_mult_29s_25s_0_7_8), .S0(s_mult_29s_25s_0_7_17), .S1(s_mult_29s_25s_0_7_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_9 (.A0(s_mult_29s_25s_0_0_19), .A1(s_mult_29s_25s_0_0_20), 
           .B0(s_mult_29s_25s_0_1_19), .B1(s_mult_29s_25s_0_1_20), .CI(co_mult_29s_25s_0_7_8), 
           .COUT(co_mult_29s_25s_0_7_9), .S0(s_mult_29s_25s_0_7_19), .S1(s_mult_29s_25s_0_7_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_10 (.A0(s_mult_29s_25s_0_0_21), .A1(s_mult_29s_25s_0_0_22), 
           .B0(s_mult_29s_25s_0_1_21), .B1(s_mult_29s_25s_0_1_22), .CI(co_mult_29s_25s_0_7_9), 
           .COUT(co_mult_29s_25s_0_7_10), .S0(s_mult_29s_25s_0_7_21), .S1(s_mult_29s_25s_0_7_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_11 (.A0(s_mult_29s_25s_0_0_23), .A1(s_mult_29s_25s_0_0_24), 
           .B0(s_mult_29s_25s_0_1_23), .B1(s_mult_29s_25s_0_1_24), .CI(co_mult_29s_25s_0_7_10), 
           .COUT(co_mult_29s_25s_0_7_11), .S0(s_mult_29s_25s_0_7_23), .S1(s_mult_29s_25s_0_7_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_12 (.A0(s_mult_29s_25s_0_0_25), .A1(s_mult_29s_25s_0_0_26), 
           .B0(s_mult_29s_25s_0_1_25), .B1(s_mult_29s_25s_0_1_26), .CI(co_mult_29s_25s_0_7_11), 
           .COUT(co_mult_29s_25s_0_7_12), .S0(s_mult_29s_25s_0_7_25), .S1(s_mult_29s_25s_0_7_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_13 (.A0(s_mult_29s_25s_0_0_27), .A1(s_mult_29s_25s_0_0_28), 
           .B0(s_mult_29s_25s_0_1_27), .B1(s_mult_29s_25s_0_1_28), .CI(co_mult_29s_25s_0_7_12), 
           .S0(s_mult_29s_25s_0_7_27), .S1(s_mult_29s_25s_0_7_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_8_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_2_12), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_6_12), .CI(GND_net), .COUT(co_mult_29s_25s_0_8_1), 
           .S1(s_mult_29s_25s_0_8_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_2 (.A0(s_mult_29s_25s_0_2_13), .A1(s_mult_29s_25s_0_2_14), 
           .B0(mult_29s_25s_0_pp_6_13), .B1(s_mult_29s_25s_0_3_14), .CI(co_mult_29s_25s_0_8_1), 
           .COUT(co_mult_29s_25s_0_8_2), .S0(s_mult_29s_25s_0_8_13), .S1(s_mult_29s_25s_0_8_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_3 (.A0(s_mult_29s_25s_0_2_15), .A1(s_mult_29s_25s_0_2_16), 
           .B0(s_mult_29s_25s_0_3_15), .B1(s_mult_29s_25s_0_3_16), .CI(co_mult_29s_25s_0_8_2), 
           .COUT(co_mult_29s_25s_0_8_3), .S0(s_mult_29s_25s_0_8_15), .S1(s_mult_29s_25s_0_8_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_4 (.A0(s_mult_29s_25s_0_2_17), .A1(s_mult_29s_25s_0_2_18), 
           .B0(s_mult_29s_25s_0_3_17), .B1(s_mult_29s_25s_0_3_18), .CI(co_mult_29s_25s_0_8_3), 
           .COUT(co_mult_29s_25s_0_8_4), .S0(s_mult_29s_25s_0_8_17), .S1(s_mult_29s_25s_0_8_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_5 (.A0(s_mult_29s_25s_0_2_19), .A1(s_mult_29s_25s_0_2_20), 
           .B0(s_mult_29s_25s_0_3_19), .B1(s_mult_29s_25s_0_3_20), .CI(co_mult_29s_25s_0_8_4), 
           .COUT(co_mult_29s_25s_0_8_5), .S0(s_mult_29s_25s_0_8_19), .S1(s_mult_29s_25s_0_8_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_6 (.A0(s_mult_29s_25s_0_2_21), .A1(s_mult_29s_25s_0_2_22), 
           .B0(s_mult_29s_25s_0_3_21), .B1(s_mult_29s_25s_0_3_22), .CI(co_mult_29s_25s_0_8_5), 
           .COUT(co_mult_29s_25s_0_8_6), .S0(s_mult_29s_25s_0_8_21), .S1(s_mult_29s_25s_0_8_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_7 (.A0(s_mult_29s_25s_0_2_23), .A1(s_mult_29s_25s_0_2_24), 
           .B0(s_mult_29s_25s_0_3_23), .B1(s_mult_29s_25s_0_3_24), .CI(co_mult_29s_25s_0_8_6), 
           .COUT(co_mult_29s_25s_0_8_7), .S0(s_mult_29s_25s_0_8_23), .S1(s_mult_29s_25s_0_8_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_8 (.A0(s_mult_29s_25s_0_2_25), .A1(s_mult_29s_25s_0_2_26), 
           .B0(s_mult_29s_25s_0_3_25), .B1(s_mult_29s_25s_0_3_26), .CI(co_mult_29s_25s_0_8_7), 
           .COUT(co_mult_29s_25s_0_8_8), .S0(s_mult_29s_25s_0_8_25), .S1(s_mult_29s_25s_0_8_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_9 (.A0(s_mult_29s_25s_0_2_27), .A1(s_mult_29s_25s_0_2_28), 
           .B0(s_mult_29s_25s_0_3_27), .B1(s_mult_29s_25s_0_3_28), .CI(co_mult_29s_25s_0_8_8), 
           .S0(s_mult_29s_25s_0_8_27), .S1(s_mult_29s_25s_0_8_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_9_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_4_20), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_10_20), .CI(GND_net), .COUT(co_mult_29s_25s_0_9_1), 
           .S1(s_mult_29s_25s_0_9_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_2 (.A0(s_mult_29s_25s_0_4_21), .A1(s_mult_29s_25s_0_4_22), 
           .B0(mult_29s_25s_0_pp_10_21), .B1(s_mult_29s_25s_0_5_22), .CI(co_mult_29s_25s_0_9_1), 
           .COUT(co_mult_29s_25s_0_9_2), .S0(s_mult_29s_25s_0_9_21), .S1(s_mult_29s_25s_0_9_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_3 (.A0(s_mult_29s_25s_0_4_23), .A1(s_mult_29s_25s_0_4_24), 
           .B0(s_mult_29s_25s_0_5_23), .B1(s_mult_29s_25s_0_5_24), .CI(co_mult_29s_25s_0_9_2), 
           .COUT(co_mult_29s_25s_0_9_3), .S0(s_mult_29s_25s_0_9_23), .S1(s_mult_29s_25s_0_9_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_4 (.A0(s_mult_29s_25s_0_4_25), .A1(s_mult_29s_25s_0_4_26), 
           .B0(s_mult_29s_25s_0_5_25), .B1(s_mult_29s_25s_0_5_26), .CI(co_mult_29s_25s_0_9_3), 
           .COUT(co_mult_29s_25s_0_9_4), .S0(s_mult_29s_25s_0_9_25), .S1(s_mult_29s_25s_0_9_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_5 (.A0(s_mult_29s_25s_0_4_27), .A1(s_mult_29s_25s_0_4_28), 
           .B0(s_mult_29s_25s_0_5_27), .B1(s_mult_29s_25s_0_5_28), .CI(co_mult_29s_25s_0_9_4), 
           .S0(s_mult_29s_25s_0_9_27), .S1(s_mult_29s_25s_0_9_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_10_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_7_8), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_4_8), .CI(GND_net), .COUT(co_mult_29s_25s_0_10_1), 
           .S1(multOut_28__N_1178[8])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_2 (.A0(s_mult_29s_25s_0_7_9), .A1(s_mult_29s_25s_0_7_10), 
           .B0(mult_29s_25s_0_pp_4_9), .B1(s_mult_29s_25s_0_2_10), .CI(co_mult_29s_25s_0_10_1), 
           .COUT(co_mult_29s_25s_0_10_2), .S0(multOut_28__N_1178[9]), .S1(multOut_28__N_1178[10])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_3 (.A0(s_mult_29s_25s_0_7_11), .A1(s_mult_29s_25s_0_7_12), 
           .B0(s_mult_29s_25s_0_2_11), .B1(s_mult_29s_25s_0_8_12), .CI(co_mult_29s_25s_0_10_2), 
           .COUT(co_mult_29s_25s_0_10_3), .S0(multOut_28__N_1178[11]), .S1(multOut_28__N_1178[12])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_4 (.A0(s_mult_29s_25s_0_7_13), .A1(s_mult_29s_25s_0_7_14), 
           .B0(s_mult_29s_25s_0_8_13), .B1(s_mult_29s_25s_0_8_14), .CI(co_mult_29s_25s_0_10_3), 
           .COUT(co_mult_29s_25s_0_10_4), .S0(multOut_28__N_1178[13]), .S1(multOut_28__N_1178[14])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_5 (.A0(s_mult_29s_25s_0_7_15), .A1(s_mult_29s_25s_0_7_16), 
           .B0(s_mult_29s_25s_0_8_15), .B1(s_mult_29s_25s_0_8_16), .CI(co_mult_29s_25s_0_10_4), 
           .COUT(co_mult_29s_25s_0_10_5), .S0(multOut_28__N_1178[15]), .S1(s_mult_29s_25s_0_10_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_6 (.A0(s_mult_29s_25s_0_7_17), .A1(s_mult_29s_25s_0_7_18), 
           .B0(s_mult_29s_25s_0_8_17), .B1(s_mult_29s_25s_0_8_18), .CI(co_mult_29s_25s_0_10_5), 
           .COUT(co_mult_29s_25s_0_10_6), .S0(s_mult_29s_25s_0_10_17), .S1(s_mult_29s_25s_0_10_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_7 (.A0(s_mult_29s_25s_0_7_19), .A1(s_mult_29s_25s_0_7_20), 
           .B0(s_mult_29s_25s_0_8_19), .B1(s_mult_29s_25s_0_8_20), .CI(co_mult_29s_25s_0_10_6), 
           .COUT(co_mult_29s_25s_0_10_7), .S0(s_mult_29s_25s_0_10_19), .S1(s_mult_29s_25s_0_10_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_8 (.A0(s_mult_29s_25s_0_7_21), .A1(s_mult_29s_25s_0_7_22), 
           .B0(s_mult_29s_25s_0_8_21), .B1(s_mult_29s_25s_0_8_22), .CI(co_mult_29s_25s_0_10_7), 
           .COUT(co_mult_29s_25s_0_10_8), .S0(s_mult_29s_25s_0_10_21), .S1(s_mult_29s_25s_0_10_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_9 (.A0(s_mult_29s_25s_0_7_23), .A1(s_mult_29s_25s_0_7_24), 
           .B0(s_mult_29s_25s_0_8_23), .B1(s_mult_29s_25s_0_8_24), .CI(co_mult_29s_25s_0_10_8), 
           .COUT(co_mult_29s_25s_0_10_9), .S0(s_mult_29s_25s_0_10_23), .S1(s_mult_29s_25s_0_10_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_10 (.A0(s_mult_29s_25s_0_7_25), .A1(s_mult_29s_25s_0_7_26), 
           .B0(s_mult_29s_25s_0_8_25), .B1(s_mult_29s_25s_0_8_26), .CI(co_mult_29s_25s_0_10_9), 
           .COUT(co_mult_29s_25s_0_10_10), .S0(s_mult_29s_25s_0_10_25), 
           .S1(s_mult_29s_25s_0_10_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_11 (.A0(s_mult_29s_25s_0_7_27), .A1(s_mult_29s_25s_0_7_28), 
           .B0(s_mult_29s_25s_0_8_27), .B1(s_mult_29s_25s_0_8_28), .CI(co_mult_29s_25s_0_10_10), 
           .S0(s_mult_29s_25s_0_10_27), .S1(s_mult_29s_25s_0_10_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_11_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_9_24), 
           .B0(GND_net), .B1(s_mult_29s_25s_0_6_24), .CI(GND_net), .COUT(co_mult_29s_25s_0_11_1), 
           .S1(s_mult_29s_25s_0_11_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_2 (.A0(s_mult_29s_25s_0_9_25), .A1(s_mult_29s_25s_0_9_26), 
           .B0(s_mult_29s_25s_0_6_25), .B1(s_mult_29s_25s_0_6_26), .CI(co_mult_29s_25s_0_11_1), 
           .COUT(co_mult_29s_25s_0_11_2), .S0(s_mult_29s_25s_0_11_25), .S1(s_mult_29s_25s_0_11_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_3 (.A0(s_mult_29s_25s_0_9_27), .A1(s_mult_29s_25s_0_9_28), 
           .B0(s_mult_29s_25s_0_6_27), .B1(s_mult_29s_25s_0_6_28), .CI(co_mult_29s_25s_0_11_2), 
           .S0(s_mult_29s_25s_0_11_27), .S1(s_mult_29s_25s_0_11_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_139_i28_3_lut (.A(n648[27]), .B(intgOut0[27]), .C(n21551), 
         .Z(n678[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i28_3_lut.init = 16'hcaca;
    LUT4 mux_135_i28_4_lut (.A(backOut2[27]), .B(backOut3[27]), .C(n21524), 
         .D(n15859), .Z(n558[27])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i28_4_lut.init = 16'hca0a;
    LUT4 mux_139_i9_3_lut (.A(n648[8]), .B(intgOut0[8]), .C(n21551), .Z(n678[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i9_3_lut.init = 16'hcaca;
    LUT4 mux_135_i9_4_lut (.A(backOut2[8]), .B(backOut3[8]), .C(n21524), 
         .D(n15859), .Z(n558[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i9_4_lut.init = 16'hca0a;
    LUT4 mux_139_i19_3_lut (.A(n648[18]), .B(intgOut0[18]), .C(n21551), 
         .Z(n678[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i19_3_lut.init = 16'hcaca;
    FADD2B Cadd_t_mult_29s_25s_0_12_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_10_16), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_8_16), .CI(GND_net), .COUT(co_t_mult_29s_25s_0_12_1), 
           .S1(multOut_28__N_1178[16])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_2 (.A0(s_mult_29s_25s_0_10_17), .A1(s_mult_29s_25s_0_10_18), 
           .B0(mult_29s_25s_0_pp_8_17), .B1(s_mult_29s_25s_0_4_18), .CI(co_t_mult_29s_25s_0_12_1), 
           .COUT(co_t_mult_29s_25s_0_12_2), .S0(multOut_28__N_1178[17]), 
           .S1(multOut_28__N_1178[18])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_3 (.A0(s_mult_29s_25s_0_10_19), .A1(s_mult_29s_25s_0_10_20), 
           .B0(s_mult_29s_25s_0_4_19), .B1(s_mult_29s_25s_0_9_20), .CI(co_t_mult_29s_25s_0_12_2), 
           .COUT(co_t_mult_29s_25s_0_12_3), .S0(multOut_28__N_1178[19]), 
           .S1(multOut_28__N_1178[20])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_4 (.A0(s_mult_29s_25s_0_10_21), .A1(s_mult_29s_25s_0_10_22), 
           .B0(s_mult_29s_25s_0_9_21), .B1(s_mult_29s_25s_0_9_22), .CI(co_t_mult_29s_25s_0_12_3), 
           .COUT(co_t_mult_29s_25s_0_12_4), .S0(multOut_28__N_1178[21]), 
           .S1(multOut_28__N_1178[22])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_5 (.A0(s_mult_29s_25s_0_10_23), .A1(s_mult_29s_25s_0_10_24), 
           .B0(s_mult_29s_25s_0_9_23), .B1(s_mult_29s_25s_0_11_24), .CI(co_t_mult_29s_25s_0_12_4), 
           .COUT(co_t_mult_29s_25s_0_12_5), .S0(multOut_28__N_1178[23]), 
           .S1(multOut_28__N_1178[24])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_6 (.A0(s_mult_29s_25s_0_10_25), .A1(s_mult_29s_25s_0_10_26), 
           .B0(s_mult_29s_25s_0_11_25), .B1(s_mult_29s_25s_0_11_26), .CI(co_t_mult_29s_25s_0_12_5), 
           .COUT(co_t_mult_29s_25s_0_12_6), .S0(multOut_28__N_1178[25]), 
           .S1(multOut_28__N_1178[26])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_7 (.A0(s_mult_29s_25s_0_10_27), .A1(s_mult_29s_25s_0_10_28), 
           .B0(s_mult_29s_25s_0_11_27), .B1(s_mult_29s_25s_0_11_28), .CI(co_t_mult_29s_25s_0_12_6), 
           .S0(multOut_28__N_1178[27]), .S1(multOut_28__N_1178[28])) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_135_i19_4_lut (.A(backOut2[18]), .B(backOut3[18]), .C(n21524), 
         .D(n15859), .Z(n558[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i19_4_lut.init = 16'hca0a;
    LUT4 mux_139_i27_3_lut (.A(n648[26]), .B(intgOut0[26]), .C(n21551), 
         .Z(n678[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i27_3_lut.init = 16'hcaca;
    LUT4 mux_135_i27_4_lut (.A(backOut2[26]), .B(backOut3[26]), .C(n21524), 
         .D(n15859), .Z(n558[26])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i27_4_lut.init = 16'hca0a;
    LUT4 mux_139_i8_3_lut (.A(n648[7]), .B(intgOut0[7]), .C(n21551), .Z(n678[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i8_3_lut.init = 16'hcaca;
    LUT4 mux_135_i8_4_lut (.A(backOut2[7]), .B(backOut3[7]), .C(n21524), 
         .D(n15859), .Z(n558[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i8_4_lut.init = 16'hca0a;
    MULT2 mult_29s_25s_0_mult_0_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_0), .CO(mco), .P0(multOut_28__N_1178[1]), 
          .P1(mult_29s_25s_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco), .CO(mco_1), .P0(mult_29s_25s_0_pp_0_3), 
          .P1(mult_29s_25s_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_1), .CO(mco_2), .P0(mult_29s_25s_0_pp_0_5), 
          .P1(mult_29s_25s_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_2), .CO(mco_3), .P0(mult_29s_25s_0_pp_0_7), 
          .P1(mult_29s_25s_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_3), .CO(mco_4), .P0(mult_29s_25s_0_pp_0_9), 
          .P1(mult_29s_25s_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_4), .CO(mco_5), .P0(mult_29s_25s_0_pp_0_11), 
          .P1(mult_29s_25s_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_5), .CO(mco_6), .P0(mult_29s_25s_0_pp_0_13), 
          .P1(mult_29s_25s_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_6), .CO(mco_7), .P0(mult_29s_25s_0_pp_0_15), 
          .P1(mult_29s_25s_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_7), .CO(mco_8), .P0(mult_29s_25s_0_pp_0_17), 
          .P1(mult_29s_25s_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_8), .CO(mco_9), .P0(mult_29s_25s_0_pp_0_19), 
          .P1(mult_29s_25s_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_9), .CO(mco_10), .P0(mult_29s_25s_0_pp_0_21), 
          .P1(mult_29s_25s_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_10), .CO(mco_11), .P0(mult_29s_25s_0_pp_0_23), 
          .P1(mult_29s_25s_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_11), .CO(mco_12), .P0(mult_29s_25s_0_pp_0_25), 
          .P1(mult_29s_25s_0_pp_0_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_13 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_12), .P0(mult_29s_25s_0_pp_0_27), .P1(mult_29s_25s_0_pp_0_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_2), .CO(mco_14), 
          .P0(mult_29s_25s_0_pp_1_3), .P1(mult_29s_25s_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_14), .CO(mco_15), .P0(mult_29s_25s_0_pp_1_5), 
          .P1(mult_29s_25s_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_15), .CO(mco_16), .P0(mult_29s_25s_0_pp_1_7), 
          .P1(mult_29s_25s_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_16), .CO(mco_17), .P0(mult_29s_25s_0_pp_1_9), 
          .P1(mult_29s_25s_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_17), .CO(mco_18), .P0(mult_29s_25s_0_pp_1_11), 
          .P1(mult_29s_25s_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_18), .CO(mco_19), .P0(mult_29s_25s_0_pp_1_13), 
          .P1(mult_29s_25s_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_19), .CO(mco_20), .P0(mult_29s_25s_0_pp_1_15), 
          .P1(mult_29s_25s_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_20), .CO(mco_21), .P0(mult_29s_25s_0_pp_1_17), 
          .P1(mult_29s_25s_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_21), .CO(mco_22), .P0(mult_29s_25s_0_pp_1_19), 
          .P1(mult_29s_25s_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_22), .CO(mco_23), .P0(mult_29s_25s_0_pp_1_21), 
          .P1(mult_29s_25s_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_23), .CO(mco_24), .P0(mult_29s_25s_0_pp_1_23), 
          .P1(mult_29s_25s_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_24), .CO(mco_25), .P0(mult_29s_25s_0_pp_1_25), 
          .P1(mult_29s_25s_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(multIn2[4]), .B2(multIn2[3]), 
          .B3(multIn2[4]), .CI(mco_25), .P0(mult_29s_25s_0_pp_1_27), .P1(mult_29s_25s_0_pp_1_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_4), .CO(mco_28), 
          .P0(mult_29s_25s_0_pp_2_5), .P1(mult_29s_25s_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_28), .CO(mco_29), .P0(mult_29s_25s_0_pp_2_7), 
          .P1(mult_29s_25s_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_29), .CO(mco_30), .P0(mult_29s_25s_0_pp_2_9), 
          .P1(mult_29s_25s_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_30), .CO(mco_31), .P0(mult_29s_25s_0_pp_2_11), 
          .P1(mult_29s_25s_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_31), .CO(mco_32), .P0(mult_29s_25s_0_pp_2_13), 
          .P1(mult_29s_25s_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_32), .CO(mco_33), .P0(mult_29s_25s_0_pp_2_15), 
          .P1(mult_29s_25s_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_33), .CO(mco_34), .P0(mult_29s_25s_0_pp_2_17), 
          .P1(mult_29s_25s_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_34), .CO(mco_35), .P0(mult_29s_25s_0_pp_2_19), 
          .P1(mult_29s_25s_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_35), .CO(mco_36), .P0(mult_29s_25s_0_pp_2_21), 
          .P1(mult_29s_25s_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_36), .CO(mco_37), .P0(mult_29s_25s_0_pp_2_23), 
          .P1(mult_29s_25s_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_37), .CO(mco_38), .P0(mult_29s_25s_0_pp_2_25), 
          .P1(mult_29s_25s_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[5]), .B1(multIn2[4]), .B2(multIn2[5]), 
          .B3(multIn2[4]), .CI(mco_38), .P0(mult_29s_25s_0_pp_2_27), .P1(mult_29s_25s_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mult_29s_25s_0_cin_lr_6), .CO(mco_42), 
          .P0(mult_29s_25s_0_pp_3_7), .P1(mult_29s_25s_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_42), .CO(mco_43), .P0(mult_29s_25s_0_pp_3_9), 
          .P1(mult_29s_25s_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_43), .CO(mco_44), .P0(mult_29s_25s_0_pp_3_11), 
          .P1(mult_29s_25s_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_44), .CO(mco_45), .P0(mult_29s_25s_0_pp_3_13), 
          .P1(mult_29s_25s_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_45), .CO(mco_46), .P0(mult_29s_25s_0_pp_3_15), 
          .P1(mult_29s_25s_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_46), .CO(mco_47), .P0(mult_29s_25s_0_pp_3_17), 
          .P1(mult_29s_25s_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_47), .CO(mco_48), .P0(mult_29s_25s_0_pp_3_19), 
          .P1(mult_29s_25s_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_48), .CO(mco_49), .P0(mult_29s_25s_0_pp_3_21), 
          .P1(mult_29s_25s_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_49), .CO(mco_50), .P0(mult_29s_25s_0_pp_3_23), 
          .P1(mult_29s_25s_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_50), .CO(mco_51), .P0(mult_29s_25s_0_pp_3_25), 
          .P1(mult_29s_25s_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_51), .P0(mult_29s_25s_0_pp_3_27), .P1(mult_29s_25s_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mult_29s_25s_0_cin_lr_8), .CO(mco_56), 
          .P0(mult_29s_25s_0_pp_4_9), .P1(mult_29s_25s_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_56), .CO(mco_57), .P0(mult_29s_25s_0_pp_4_11), 
          .P1(mult_29s_25s_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_57), .CO(mco_58), .P0(mult_29s_25s_0_pp_4_13), 
          .P1(mult_29s_25s_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_58), .CO(mco_59), .P0(mult_29s_25s_0_pp_4_15), 
          .P1(mult_29s_25s_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_59), .CO(mco_60), .P0(mult_29s_25s_0_pp_4_17), 
          .P1(mult_29s_25s_0_pp_4_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_60), .CO(mco_61), .P0(mult_29s_25s_0_pp_4_19), 
          .P1(mult_29s_25s_0_pp_4_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_61), .CO(mco_62), .P0(mult_29s_25s_0_pp_4_21), 
          .P1(mult_29s_25s_0_pp_4_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_62), .CO(mco_63), .P0(mult_29s_25s_0_pp_4_23), 
          .P1(mult_29s_25s_0_pp_4_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_63), .CO(mco_64), .P0(mult_29s_25s_0_pp_4_25), 
          .P1(mult_29s_25s_0_pp_4_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[4]), .B1(multIn2[6]), .B2(multIn2[4]), 
          .B3(multIn2[6]), .CI(mco_64), .P0(mult_29s_25s_0_pp_4_27), .P1(mult_29s_25s_0_pp_4_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 i10352_3_lut_4_lut (.A(n1187[15]), .B(n30), .C(n18815), .D(clk_N_683_enable_392), 
         .Z(n12655)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(342[7:42])
    defparam i10352_3_lut_4_lut.init = 16'hf700;
    MULT2 mult_29s_25s_0_mult_10_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_10), .CO(mco_70), .P0(mult_29s_25s_0_pp_5_11), 
          .P1(mult_29s_25s_0_pp_5_12)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_70), .CO(mco_71), .P0(mult_29s_25s_0_pp_5_13), 
          .P1(mult_29s_25s_0_pp_5_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_71), .CO(mco_72), .P0(mult_29s_25s_0_pp_5_15), 
          .P1(mult_29s_25s_0_pp_5_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_72), .CO(mco_73), .P0(mult_29s_25s_0_pp_5_17), 
          .P1(mult_29s_25s_0_pp_5_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_73), .CO(mco_74), .P0(mult_29s_25s_0_pp_5_19), 
          .P1(mult_29s_25s_0_pp_5_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_74), .CO(mco_75), .P0(mult_29s_25s_0_pp_5_21), 
          .P1(mult_29s_25s_0_pp_5_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_75), .CO(mco_76), .P0(mult_29s_25s_0_pp_5_23), 
          .P1(mult_29s_25s_0_pp_5_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_76), .CO(mco_77), .P0(mult_29s_25s_0_pp_5_25), 
          .P1(mult_29s_25s_0_pp_5_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[6]), .B1(GND_net), .B2(multIn2[6]), 
          .B3(GND_net), .CI(mco_77), .P0(mult_29s_25s_0_pp_5_27), .P1(mult_29s_25s_0_pp_5_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_139_i18_3_lut (.A(n648[17]), .B(intgOut0[17]), .C(n21551), 
         .Z(n678[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i18_3_lut.init = 16'hcaca;
    MULT2 mult_29s_25s_0_mult_12_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_12), .CO(mco_84), .P0(mult_29s_25s_0_pp_6_13), 
          .P1(mult_29s_25s_0_pp_6_14)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_84), .CO(mco_85), .P0(mult_29s_25s_0_pp_6_15), 
          .P1(mult_29s_25s_0_pp_6_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_85), .CO(mco_86), .P0(mult_29s_25s_0_pp_6_17), 
          .P1(mult_29s_25s_0_pp_6_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_86), .CO(mco_87), .P0(mult_29s_25s_0_pp_6_19), 
          .P1(mult_29s_25s_0_pp_6_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_87), .CO(mco_88), .P0(mult_29s_25s_0_pp_6_21), 
          .P1(mult_29s_25s_0_pp_6_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_88), .CO(mco_89), .P0(mult_29s_25s_0_pp_6_23), 
          .P1(mult_29s_25s_0_pp_6_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_89), .CO(mco_90), .P0(mult_29s_25s_0_pp_6_25), 
          .P1(mult_29s_25s_0_pp_6_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_90), .P0(mult_29s_25s_0_pp_6_27), .P1(mult_29s_25s_0_pp_6_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_135_i18_4_lut (.A(backOut2[17]), .B(backOut3[17]), .C(n21524), 
         .D(n15859), .Z(n558[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i18_4_lut.init = 16'hca0a;
    MULT2 mult_29s_25s_0_mult_14_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_14), .CO(mco_98), .P0(mult_29s_25s_0_pp_7_15), 
          .P1(mult_29s_25s_0_pp_7_16)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_98), .CO(mco_99), .P0(mult_29s_25s_0_pp_7_17), 
          .P1(mult_29s_25s_0_pp_7_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_99), .CO(mco_100), .P0(mult_29s_25s_0_pp_7_19), 
          .P1(mult_29s_25s_0_pp_7_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_100), .CO(mco_101), .P0(mult_29s_25s_0_pp_7_21), 
          .P1(mult_29s_25s_0_pp_7_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_101), .CO(mco_102), .P0(mult_29s_25s_0_pp_7_23), 
          .P1(mult_29s_25s_0_pp_7_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_102), .CO(mco_103), .P0(mult_29s_25s_0_pp_7_25), 
          .P1(mult_29s_25s_0_pp_7_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_103), .P0(mult_29s_25s_0_pp_7_27), .P1(mult_29s_25s_0_pp_7_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 i13925_4_lut_4_lut (.A(n920), .B(n3635), .C(addOut[14]), .D(n22208), 
         .Z(intgOut0_28__N_735[14])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13925_4_lut_4_lut.init = 16'h00ba;
    MULT2 mult_29s_25s_0_mult_16_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_16), .CO(mco_112), .P0(mult_29s_25s_0_pp_8_17), 
          .P1(mult_29s_25s_0_pp_8_18)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_112), .CO(mco_113), .P0(mult_29s_25s_0_pp_8_19), 
          .P1(mult_29s_25s_0_pp_8_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_113), .CO(mco_114), .P0(mult_29s_25s_0_pp_8_21), 
          .P1(mult_29s_25s_0_pp_8_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_114), .CO(mco_115), .P0(mult_29s_25s_0_pp_8_23), 
          .P1(mult_29s_25s_0_pp_8_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_115), .CO(mco_116), .P0(mult_29s_25s_0_pp_8_25), 
          .P1(mult_29s_25s_0_pp_8_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_116), .P0(mult_29s_25s_0_pp_8_27), .P1(mult_29s_25s_0_pp_8_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_139_i26_3_lut (.A(n648[25]), .B(intgOut0[25]), .C(n21551), 
         .Z(n678[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i26_3_lut.init = 16'hcaca;
    LUT4 mux_135_i26_4_lut (.A(backOut2[25]), .B(backOut3[25]), .C(n21524), 
         .D(n15859), .Z(n558[25])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i26_4_lut.init = 16'hca0a;
    MULT2 mult_29s_25s_0_mult_18_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_18), .CO(mco_126), .P0(mult_29s_25s_0_pp_9_19), 
          .P1(mult_29s_25s_0_pp_9_20)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_126), .CO(mco_127), .P0(mult_29s_25s_0_pp_9_21), 
          .P1(mult_29s_25s_0_pp_9_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_127), .CO(mco_128), .P0(mult_29s_25s_0_pp_9_23), 
          .P1(mult_29s_25s_0_pp_9_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_128), .CO(mco_129), .P0(mult_29s_25s_0_pp_9_25), 
          .P1(mult_29s_25s_0_pp_9_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_129), .P0(mult_29s_25s_0_pp_9_27), .P1(mult_29s_25s_0_pp_9_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_139_i7_3_lut (.A(n648[6]), .B(intgOut0[6]), .C(n21551), .Z(n678[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i7_3_lut.init = 16'hcaca;
    MULT2 mult_29s_25s_0_mult_20_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_20), .CO(mco_140), .P0(mult_29s_25s_0_pp_10_21), 
          .P1(mult_29s_25s_0_pp_10_22)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_140), .CO(mco_141), .P0(mult_29s_25s_0_pp_10_23), 
          .P1(mult_29s_25s_0_pp_10_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_141), .CO(mco_142), .P0(mult_29s_25s_0_pp_10_25), 
          .P1(mult_29s_25s_0_pp_10_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_142), .P0(mult_29s_25s_0_pp_10_27), .P1(mult_29s_25s_0_pp_10_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 mux_135_i7_4_lut (.A(backOut2[6]), .B(backOut3[6]), .C(n21524), 
         .D(n15859), .Z(n558[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i7_4_lut.init = 16'hca0a;
    LUT4 i17866_4_lut_4_lut (.A(n21510), .B(n20450), .C(n21526), .D(n21543), 
         .Z(n20579)) /* synthesis lut_function=(!(A (C (D))+!A !(B+!(C (D))))) */ ;
    defparam i17866_4_lut_4_lut.init = 16'h4fff;
    MULT2 mult_29s_25s_0_mult_22_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_22), .CO(mco_154), .P0(mult_29s_25s_0_pp_11_23), 
          .P1(mult_29s_25s_0_pp_11_24)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_154), .CO(mco_155), .P0(mult_29s_25s_0_pp_11_25), 
          .P1(mult_29s_25s_0_pp_11_26)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_155), .P0(mult_29s_25s_0_pp_11_27), .P1(mult_29s_25s_0_pp_11_28)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 i17774_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[25]), .D(n558[25]), 
         .Z(addIn2_28__N_1337[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17774_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17726_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[16]), .D(n558[16]), 
         .Z(addIn2_28__N_1337[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17726_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17752_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[2]), .D(n558[2]), 
         .Z(addIn2_28__N_1337[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17752_3_lut_4_lut.init = 16'hf1e0;
    FADD2B mult_29s_25s_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(229[14:21])
    LUT4 i17758_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[17]), .D(n558[17]), 
         .Z(addIn2_28__N_1337[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17758_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_50 (.A(n920), .B(n3635), .C(addOut[2]), 
         .D(n22208), .Z(intgOut0_28__N_735[2])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_50.init = 16'h0010;
    LUT4 mux_139_i17_3_lut (.A(n648[16]), .B(intgOut0[16]), .C(n21551), 
         .Z(n678[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i17_3_lut.init = 16'hcaca;
    LUT4 mux_135_i17_4_lut (.A(backOut2[16]), .B(backOut3[16]), .C(n21524), 
         .D(n15859), .Z(n558[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i17_4_lut.init = 16'hca0a;
    PFUMX mux_1193_i11 (.BLUT(n5109), .ALUT(n5067), .C0(n2436), .Z(n5157));
    LUT4 i17734_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[12]), .D(n558[12]), 
         .Z(addIn2_28__N_1337[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17734_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17772_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[24]), .D(n558[24]), 
         .Z(addIn2_28__N_1337[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17772_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17728_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[15]), .D(n558[15]), 
         .Z(addIn2_28__N_1337[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17728_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17754_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[6]), .D(n558[6]), 
         .Z(addIn2_28__N_1337[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17754_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_1193_i10 (.BLUT(n5107), .ALUT(n5065), .C0(n2436), .Z(n5155));
    LUT4 i17760_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[18]), .D(n558[18]), 
         .Z(addIn2_28__N_1337[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17760_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17748_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[3]), .D(n558[3]), 
         .Z(addIn2_28__N_1337[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17748_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17778_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[27]), .D(n558[27]), 
         .Z(addIn2_28__N_1337[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17778_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_1193_i9 (.BLUT(n5105), .ALUT(n5063), .C0(n2436), .Z(n5153));
    LUT4 i17780_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[28]), .D(n558[28]), 
         .Z(addIn2_28__N_1337[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17780_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i25_3_lut (.A(n648[24]), .B(intgOut0[24]), .C(n21551), 
         .Z(n678[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i25_3_lut.init = 16'hcaca;
    LUT4 i17756_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[8]), .D(n558[8]), 
         .Z(addIn2_28__N_1337[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17756_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i25_4_lut (.A(backOut2[24]), .B(backOut3[24]), .C(n21524), 
         .D(n15859), .Z(n558[24])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i25_4_lut.init = 16'hca0a;
    LUT4 i13927_4_lut_4_lut (.A(n920), .B(n3635), .C(addOut[16]), .D(n22208), 
         .Z(intgOut0_28__N_735[16])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13927_4_lut_4_lut.init = 16'h00ba;
    LUT4 i17736_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[11]), .D(n558[11]), 
         .Z(addIn2_28__N_1337[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17736_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX addOut_2063__i0 (.D(n121[0]), .CK(clk_N_683), .Q(addOut[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i0.GSR = "ENABLED";
    LUT4 i17766_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[21]), .D(n558[21]), 
         .Z(addIn2_28__N_1337[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17766_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_1193_i8 (.BLUT(n5103), .ALUT(n5061), .C0(n2436), .Z(n5151));
    LUT4 i17744_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[5]), .D(n558[5]), 
         .Z(addIn2_28__N_1337[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17744_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17764_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[20]), .D(n558[20]), 
         .Z(addIn2_28__N_1337[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17764_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i6_3_lut (.A(n648[5]), .B(intgOut0[5]), .C(n21551), .Z(n678[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 187[26])
    defparam mux_139_i6_3_lut.init = 16'hcaca;
    LUT4 i17730_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[14]), .D(n558[14]), 
         .Z(addIn2_28__N_1337[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17730_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17776_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[26]), .D(n558[26]), 
         .Z(addIn2_28__N_1337[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17776_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_51 (.A(n920), .B(n3635), .C(addOut[3]), 
         .D(n22208), .Z(intgOut0_28__N_735[3])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_51.init = 16'h0010;
    LUT4 i17724_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[0]), .D(n558[0]), 
         .Z(addIn2_28__N_1337[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17724_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17738_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[10]), .D(n558[10]), 
         .Z(addIn2_28__N_1337[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17738_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_1193_i7 (.BLUT(n5101), .ALUT(n5059), .C0(n2436), .Z(n5149));
    LUT4 i17762_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[19]), .D(n558[19]), 
         .Z(addIn2_28__N_1337[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17762_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17750_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[7]), .D(n558[7]), 
         .Z(addIn2_28__N_1337[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17750_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17770_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[23]), .D(n558[23]), 
         .Z(addIn2_28__N_1337[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17770_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17742_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[1]), .D(n558[1]), 
         .Z(addIn2_28__N_1337[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17742_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17740_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[9]), .D(n558[9]), 
         .Z(addIn2_28__N_1337[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17740_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i6_4_lut (.A(backOut2[5]), .B(backOut3[5]), .C(n21524), 
         .D(n15859), .Z(n558[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 191[27])
    defparam mux_135_i6_4_lut.init = 16'hca0a;
    PFUMX mux_1193_i6 (.BLUT(n5099), .ALUT(n5057), .C0(n2436), .Z(n5147));
    LUT4 i17746_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[4]), .D(n558[4]), 
         .Z(addIn2_28__N_1337[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17746_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17768_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[22]), .D(n558[22]), 
         .Z(addIn2_28__N_1337[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17768_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17732_3_lut_4_lut (.A(n21551), .B(n21520), .C(n678[13]), .D(n558[13]), 
         .Z(addIn2_28__N_1337[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(184[17] 186[26])
    defparam i17732_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_1193_i5 (.BLUT(n5097), .ALUT(n5055), .C0(n2436), .Z(n5145));
    LUT4 i13928_4_lut_4_lut (.A(n920), .B(n3635), .C(addOut[17]), .D(n22208), 
         .Z(intgOut0_28__N_735[17])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13928_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_1188_i11_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m4[10]), .Z(n5109)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i11_3_lut_4_lut.init = 16'hf780;
    FD1P3AX backOut0_i0_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_73), 
            .CK(clk_N_683), .Q(backOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut0_i0_i1.GSR = "DISABLED";
    FD1S3AX multOut_i1 (.D(multOut_28__N_1178[1]), .CK(clk_N_683), .Q(multOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(n920), .B(n3635), .C(addOut[4]), 
         .D(n22208), .Z(intgOut0_28__N_735[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'h0010;
    LUT4 mux_1799_i1_4_lut (.A(\speed_m4[0] ), .B(\speed_m3[0] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i1_4_lut.init = 16'hcac0;
    LUT4 mux_1799_i4_3_lut (.A(\speed_m3[3] ), .B(\speed_m2[3] ), .C(n4138), 
         .Z(subIn2_24__N_1301[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i4_3_lut.init = 16'hcaca;
    LUT4 i13929_4_lut_4_lut (.A(n920), .B(n3635), .C(addOut[18]), .D(n22208), 
         .Z(intgOut0_28__N_735[18])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13929_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_1798_i13_3_lut_4_lut_4_lut (.A(n21508), .B(\speed_m4[12] ), 
         .C(n4132), .D(n21510), .Z(n3690[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam mux_1798_i13_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_1799_i8_3_lut (.A(\speed_m3[7] ), .B(\speed_m2[7] ), .C(n4138), 
         .Z(subIn2_24__N_1301[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1799_i9_3_lut (.A(\speed_m3[8] ), .B(\speed_m2[8] ), .C(n4138), 
         .Z(subIn2_24__N_1301[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1799_i10_3_lut (.A(\speed_m3[9] ), .B(\speed_m2[9] ), .C(n4138), 
         .Z(subIn2_24__N_1301[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1799_i13_3_lut (.A(\speed_m3[12] ), .B(\speed_m2[12] ), .C(n4138), 
         .Z(subIn2_24__N_1301[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1798_i10_3_lut_4_lut_4_lut (.A(n21508), .B(\speed_m4[9] ), 
         .C(n4132), .D(n21510), .Z(n3690[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam mux_1798_i10_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_1798_i9_3_lut_4_lut_4_lut (.A(n21508), .B(\speed_m4[8] ), .C(n4132), 
         .D(n21510), .Z(n3690[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam mux_1798_i9_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_1799_i19_4_lut (.A(\speed_m4[18] ), .B(\speed_m3[18] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i19_4_lut.init = 16'hcac0;
    LUT4 mux_1798_i8_3_lut_4_lut_4_lut (.A(n21508), .B(\speed_m4[7] ), .C(n4132), 
         .D(n21510), .Z(n3690[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam mux_1798_i8_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_1798_i4_3_lut_4_lut_4_lut (.A(n21508), .B(\speed_m4[3] ), .C(n4132), 
         .D(n21510), .Z(n3690[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam mux_1798_i4_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i7_4_lut_adj_53 (.A(Out0[3]), .B(n14_adj_1830), .C(n10_adj_1831), 
         .D(Out0[4]), .Z(n18864)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam i7_4_lut_adj_53.init = 16'hfffe;
    LUT4 mux_1799_i18_4_lut (.A(\speed_m4[17] ), .B(\speed_m3[17] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i18_4_lut.init = 16'hcac0;
    LUT4 i6_4_lut_adj_54 (.A(Out0[11]), .B(Out0[7]), .C(Out0[2]), .D(Out0[10]), 
         .Z(n14_adj_1830)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam i6_4_lut_adj_54.init = 16'hfffe;
    LUT4 i2_2_lut_adj_55 (.A(Out0[9]), .B(Out0[1]), .Z(n10_adj_1831)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam i2_2_lut_adj_55.init = 16'heeee;
    LUT4 mux_1799_i17_4_lut (.A(\speed_m4[16] ), .B(\speed_m3[16] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i17_4_lut.init = 16'hcac0;
    PFUMX mux_1193_i4 (.BLUT(n5095), .ALUT(n5053), .C0(n2436), .Z(n5143));
    LUT4 mux_1799_i16_4_lut (.A(\speed_m4[15] ), .B(\speed_m3[15] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i16_4_lut.init = 16'hcac0;
    PFUMX mux_1193_i3 (.BLUT(n5093), .ALUT(n5051), .C0(n2436), .Z(n5141));
    LUT4 i4_4_lut_adj_56 (.A(Out0[5]), .B(Out0[6]), .C(Out0[0]), .D(n6_adj_1832), 
         .Z(n18865)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam i4_4_lut_adj_56.init = 16'hfffe;
    FD1S3AX multOut_i2 (.D(multOut_28__N_1178[2]), .CK(clk_N_683), .Q(multOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i2.GSR = "ENABLED";
    FD1S3AX multOut_i3 (.D(multOut_28__N_1178[3]), .CK(clk_N_683), .Q(multOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i3.GSR = "ENABLED";
    FD1S3AX multOut_i4 (.D(multOut_28__N_1178[4]), .CK(clk_N_683), .Q(multOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i4.GSR = "ENABLED";
    FD1S3AX multOut_i5 (.D(multOut_28__N_1178[5]), .CK(clk_N_683), .Q(multOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i5.GSR = "ENABLED";
    FD1S3AX multOut_i6 (.D(multOut_28__N_1178[6]), .CK(clk_N_683), .Q(multOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i6.GSR = "ENABLED";
    FD1S3AX multOut_i7 (.D(multOut_28__N_1178[7]), .CK(clk_N_683), .Q(multOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i7.GSR = "ENABLED";
    FD1S3AX multOut_i8 (.D(multOut_28__N_1178[8]), .CK(clk_N_683), .Q(multOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i8.GSR = "ENABLED";
    FD1S3AX multOut_i9 (.D(multOut_28__N_1178[9]), .CK(clk_N_683), .Q(multOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i9.GSR = "ENABLED";
    FD1S3AX multOut_i10 (.D(multOut_28__N_1178[10]), .CK(clk_N_683), .Q(multOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i10.GSR = "ENABLED";
    FD1S3AX multOut_i11 (.D(multOut_28__N_1178[11]), .CK(clk_N_683), .Q(multOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i11.GSR = "ENABLED";
    FD1S3AX multOut_i12 (.D(multOut_28__N_1178[12]), .CK(clk_N_683), .Q(multOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i12.GSR = "ENABLED";
    FD1S3AX multOut_i13 (.D(multOut_28__N_1178[13]), .CK(clk_N_683), .Q(multOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i13.GSR = "ENABLED";
    FD1S3AX multOut_i14 (.D(multOut_28__N_1178[14]), .CK(clk_N_683), .Q(multOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i14.GSR = "ENABLED";
    FD1S3AX multOut_i15 (.D(multOut_28__N_1178[15]), .CK(clk_N_683), .Q(multOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i15.GSR = "ENABLED";
    FD1S3AX multOut_i16 (.D(multOut_28__N_1178[16]), .CK(clk_N_683), .Q(multOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i16.GSR = "ENABLED";
    FD1S3AX multOut_i17 (.D(multOut_28__N_1178[17]), .CK(clk_N_683), .Q(multOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i17.GSR = "ENABLED";
    FD1S3AX multOut_i18 (.D(multOut_28__N_1178[18]), .CK(clk_N_683), .Q(multOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i18.GSR = "ENABLED";
    FD1S3AX multOut_i19 (.D(multOut_28__N_1178[19]), .CK(clk_N_683), .Q(multOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i19.GSR = "ENABLED";
    FD1S3AX multOut_i20 (.D(multOut_28__N_1178[20]), .CK(clk_N_683), .Q(multOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i20.GSR = "ENABLED";
    FD1S3AX multOut_i21 (.D(multOut_28__N_1178[21]), .CK(clk_N_683), .Q(multOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i21.GSR = "ENABLED";
    FD1S3AX multOut_i22 (.D(multOut_28__N_1178[22]), .CK(clk_N_683), .Q(multOut[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i22.GSR = "ENABLED";
    FD1S3AX multOut_i23 (.D(multOut_28__N_1178[23]), .CK(clk_N_683), .Q(multOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i23.GSR = "ENABLED";
    FD1S3AX multOut_i24 (.D(multOut_28__N_1178[24]), .CK(clk_N_683), .Q(multOut[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i24.GSR = "ENABLED";
    FD1S3AX multOut_i25 (.D(multOut_28__N_1178[25]), .CK(clk_N_683), .Q(multOut[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i25.GSR = "ENABLED";
    FD1S3AX multOut_i26 (.D(multOut_28__N_1178[26]), .CK(clk_N_683), .Q(multOut[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i26.GSR = "ENABLED";
    FD1S3AX multOut_i27 (.D(multOut_28__N_1178[27]), .CK(clk_N_683), .Q(multOut[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i27.GSR = "ENABLED";
    FD1S3AX multOut_i28 (.D(multOut_28__N_1178[28]), .CK(clk_N_683), .Q(multOut[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam multOut_i28.GSR = "ENABLED";
    FD1P3AX intgOut0_i1 (.D(intgOut0_28__N_735[1]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i1.GSR = "ENABLED";
    FD1P3AX intgOut0_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i2.GSR = "ENABLED";
    FD1P3AX intgOut0_i3 (.D(intgOut0_28__N_735[3]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i3.GSR = "ENABLED";
    FD1P3AX intgOut0_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i4.GSR = "ENABLED";
    FD1P3AX intgOut0_i5 (.D(intgOut0_28__N_735[5]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i5.GSR = "ENABLED";
    FD1P3AX intgOut0_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i6.GSR = "ENABLED";
    FD1P3AX intgOut0_i7 (.D(intgOut0_28__N_735[7]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i7.GSR = "ENABLED";
    FD1P3AX intgOut0_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i8.GSR = "ENABLED";
    FD1P3AX intgOut0_i9 (.D(intgOut0_28__N_735[9]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i9.GSR = "ENABLED";
    FD1P3AX intgOut0_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i10.GSR = "ENABLED";
    FD1P3AX intgOut0_i11 (.D(intgOut0_28__N_735[11]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i11.GSR = "ENABLED";
    FD1P3AX intgOut0_i12 (.D(intgOut0_28__N_735[12]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i12.GSR = "ENABLED";
    FD1P3AX intgOut0_i13 (.D(intgOut0_28__N_735[13]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i13.GSR = "ENABLED";
    FD1P3AX intgOut0_i14 (.D(intgOut0_28__N_735[14]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i14.GSR = "ENABLED";
    FD1P3AX intgOut0_i15 (.D(intgOut0_28__N_735[15]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i15.GSR = "ENABLED";
    FD1P3AX intgOut0_i16 (.D(intgOut0_28__N_735[16]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i16.GSR = "ENABLED";
    FD1P3AX intgOut0_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i17.GSR = "ENABLED";
    FD1P3AX intgOut0_i18 (.D(intgOut0_28__N_735[18]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i18.GSR = "ENABLED";
    FD1P3AX intgOut0_i19 (.D(intgOut0_28__N_735[19]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i19.GSR = "ENABLED";
    FD1P3AX intgOut0_i20 (.D(intgOut0_28__N_735[20]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i20.GSR = "ENABLED";
    FD1P3AX intgOut0_i21 (.D(intgOut0_28__N_735[21]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i21.GSR = "ENABLED";
    FD1P3AX intgOut0_i22 (.D(intgOut0_28__N_735[22]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i22.GSR = "ENABLED";
    FD1P3AX intgOut0_i23 (.D(intgOut0_28__N_735[23]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i23.GSR = "ENABLED";
    FD1P3AX intgOut0_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i24.GSR = "ENABLED";
    FD1P3AX intgOut0_i25 (.D(intgOut0_28__N_735[25]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i25.GSR = "ENABLED";
    FD1P3AX intgOut0_i26 (.D(intgOut0_28__N_735[26]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i26.GSR = "ENABLED";
    FD1P3AX intgOut0_i27 (.D(intgOut0_28__N_735[27]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i27.GSR = "ENABLED";
    FD1P3AX intgOut0_i28 (.D(intgOut0_28__N_735[28]), .SP(clk_N_683_enable_101), 
            .CK(clk_N_683), .Q(intgOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut0_i28.GSR = "ENABLED";
    FD1P3AX intgOut1_i1 (.D(intgOut0_28__N_735[1]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i1.GSR = "ENABLED";
    FD1P3AX intgOut1_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i2.GSR = "ENABLED";
    FD1P3AX intgOut1_i3 (.D(intgOut0_28__N_735[3]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i3.GSR = "ENABLED";
    FD1P3AX intgOut1_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i4.GSR = "ENABLED";
    FD1P3AX intgOut1_i5 (.D(intgOut0_28__N_735[5]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i5.GSR = "ENABLED";
    FD1P3AX intgOut1_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i6.GSR = "ENABLED";
    FD1P3AX intgOut1_i7 (.D(intgOut0_28__N_735[7]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i7.GSR = "ENABLED";
    FD1P3AX intgOut1_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i8.GSR = "ENABLED";
    FD1P3AX intgOut1_i9 (.D(intgOut0_28__N_735[9]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i9.GSR = "ENABLED";
    FD1P3AX intgOut1_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i10.GSR = "ENABLED";
    FD1P3AX intgOut1_i11 (.D(intgOut0_28__N_735[11]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i11.GSR = "ENABLED";
    FD1P3AX intgOut1_i12 (.D(intgOut0_28__N_735[12]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i12.GSR = "ENABLED";
    FD1P3AX intgOut1_i13 (.D(intgOut0_28__N_735[13]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i13.GSR = "ENABLED";
    FD1P3AX intgOut1_i14 (.D(intgOut0_28__N_735[14]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i14.GSR = "ENABLED";
    FD1P3AX intgOut1_i15 (.D(intgOut0_28__N_735[15]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i15.GSR = "ENABLED";
    FD1P3AX intgOut1_i16 (.D(intgOut0_28__N_735[16]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i16.GSR = "ENABLED";
    FD1P3AX intgOut1_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i17.GSR = "ENABLED";
    FD1P3AX intgOut1_i18 (.D(intgOut0_28__N_735[18]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i18.GSR = "ENABLED";
    FD1P3AX intgOut1_i19 (.D(intgOut0_28__N_735[19]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i19.GSR = "ENABLED";
    FD1P3AX intgOut1_i20 (.D(intgOut0_28__N_735[20]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i20.GSR = "ENABLED";
    FD1P3AX intgOut1_i21 (.D(intgOut0_28__N_735[21]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i21.GSR = "ENABLED";
    FD1P3AX intgOut1_i22 (.D(intgOut0_28__N_735[22]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i22.GSR = "ENABLED";
    FD1P3AX intgOut1_i23 (.D(intgOut0_28__N_735[23]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i23.GSR = "ENABLED";
    FD1P3AX intgOut1_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i24.GSR = "ENABLED";
    FD1P3AX intgOut1_i25 (.D(intgOut0_28__N_735[25]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i25.GSR = "ENABLED";
    FD1P3AX intgOut1_i26 (.D(intgOut0_28__N_735[26]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i26.GSR = "ENABLED";
    FD1P3AX intgOut1_i27 (.D(intgOut0_28__N_735[27]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i27.GSR = "ENABLED";
    FD1P3AX intgOut1_i28 (.D(intgOut0_28__N_735[28]), .SP(clk_N_683_enable_129), 
            .CK(clk_N_683), .Q(intgOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut1_i28.GSR = "ENABLED";
    FD1P3AX intgOut2_i1 (.D(intgOut0_28__N_735[1]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i1.GSR = "ENABLED";
    FD1P3AX intgOut2_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i2.GSR = "ENABLED";
    FD1P3AX intgOut2_i3 (.D(intgOut0_28__N_735[3]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i3.GSR = "ENABLED";
    FD1P3AX intgOut2_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i4.GSR = "ENABLED";
    FD1P3AX intgOut2_i5 (.D(intgOut0_28__N_735[5]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i5.GSR = "ENABLED";
    FD1P3AX intgOut2_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i6.GSR = "ENABLED";
    FD1P3AX intgOut2_i7 (.D(intgOut0_28__N_735[7]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i7.GSR = "ENABLED";
    FD1P3AX intgOut2_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i8.GSR = "ENABLED";
    FD1P3AX intgOut2_i9 (.D(intgOut0_28__N_735[9]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i9.GSR = "ENABLED";
    FD1P3AX intgOut2_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i10.GSR = "ENABLED";
    FD1P3AX intgOut2_i11 (.D(intgOut0_28__N_735[11]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i11.GSR = "ENABLED";
    FD1P3AX intgOut2_i12 (.D(intgOut0_28__N_735[12]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i12.GSR = "ENABLED";
    FD1P3AX intgOut2_i13 (.D(intgOut0_28__N_735[13]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i13.GSR = "ENABLED";
    FD1P3AX intgOut2_i14 (.D(intgOut0_28__N_735[14]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i14.GSR = "ENABLED";
    FD1P3AX intgOut2_i15 (.D(intgOut0_28__N_735[15]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i15.GSR = "ENABLED";
    FD1P3AX intgOut2_i16 (.D(intgOut0_28__N_735[16]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i16.GSR = "ENABLED";
    FD1P3AX intgOut2_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i17.GSR = "ENABLED";
    FD1P3AX intgOut2_i18 (.D(intgOut0_28__N_735[18]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i18.GSR = "ENABLED";
    FD1P3AX intgOut2_i19 (.D(intgOut0_28__N_735[19]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i19.GSR = "ENABLED";
    FD1P3AX intgOut2_i20 (.D(intgOut0_28__N_735[20]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i20.GSR = "ENABLED";
    FD1P3AX intgOut2_i21 (.D(intgOut0_28__N_735[21]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i21.GSR = "ENABLED";
    FD1P3AX intgOut2_i22 (.D(intgOut0_28__N_735[22]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i22.GSR = "ENABLED";
    FD1P3AX intgOut2_i23 (.D(intgOut0_28__N_735[23]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i23.GSR = "ENABLED";
    FD1P3AX intgOut2_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i24.GSR = "ENABLED";
    FD1P3AX intgOut2_i25 (.D(intgOut0_28__N_735[25]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i25.GSR = "ENABLED";
    FD1P3AX intgOut2_i26 (.D(intgOut0_28__N_735[26]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i26.GSR = "ENABLED";
    FD1P3AX intgOut2_i27 (.D(intgOut0_28__N_735[27]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i27.GSR = "ENABLED";
    FD1P3AX intgOut2_i28 (.D(intgOut0_28__N_735[28]), .SP(clk_N_683_enable_157), 
            .CK(clk_N_683), .Q(intgOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut2_i28.GSR = "ENABLED";
    FD1P3AX intgOut3_i1 (.D(intgOut0_28__N_735[1]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i1.GSR = "ENABLED";
    FD1P3AX intgOut3_i2 (.D(intgOut0_28__N_735[2]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i2.GSR = "ENABLED";
    FD1P3AX intgOut3_i3 (.D(intgOut0_28__N_735[3]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i3.GSR = "ENABLED";
    FD1P3AX intgOut3_i4 (.D(intgOut0_28__N_735[4]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i4.GSR = "ENABLED";
    FD1P3AX intgOut3_i5 (.D(intgOut0_28__N_735[5]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i5.GSR = "ENABLED";
    FD1P3AX intgOut3_i6 (.D(intgOut0_28__N_735[6]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i6.GSR = "ENABLED";
    FD1P3AX intgOut3_i7 (.D(intgOut0_28__N_735[7]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i7.GSR = "ENABLED";
    FD1P3AX intgOut3_i8 (.D(intgOut0_28__N_735[8]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i8.GSR = "ENABLED";
    FD1P3AX intgOut3_i9 (.D(intgOut0_28__N_735[9]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i9.GSR = "ENABLED";
    FD1P3AX intgOut3_i10 (.D(intgOut0_28__N_735[10]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i10.GSR = "ENABLED";
    FD1P3AX intgOut3_i11 (.D(intgOut0_28__N_735[11]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i11.GSR = "ENABLED";
    FD1P3AX intgOut3_i12 (.D(intgOut0_28__N_735[12]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i12.GSR = "ENABLED";
    FD1P3AX intgOut3_i13 (.D(intgOut0_28__N_735[13]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i13.GSR = "ENABLED";
    FD1P3AX intgOut3_i14 (.D(intgOut0_28__N_735[14]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i14.GSR = "ENABLED";
    FD1P3AX intgOut3_i15 (.D(intgOut0_28__N_735[15]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i15.GSR = "ENABLED";
    FD1P3AX intgOut3_i16 (.D(intgOut0_28__N_735[16]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i16.GSR = "ENABLED";
    FD1P3AX intgOut3_i17 (.D(intgOut0_28__N_735[17]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i17.GSR = "ENABLED";
    FD1P3AX intgOut3_i18 (.D(intgOut0_28__N_735[18]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i18.GSR = "ENABLED";
    FD1P3AX intgOut3_i19 (.D(intgOut0_28__N_735[19]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i19.GSR = "ENABLED";
    FD1P3AX intgOut3_i20 (.D(intgOut0_28__N_735[20]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i20.GSR = "ENABLED";
    FD1P3AX intgOut3_i21 (.D(intgOut0_28__N_735[21]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i21.GSR = "ENABLED";
    FD1P3AX intgOut3_i22 (.D(intgOut0_28__N_735[22]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i22.GSR = "ENABLED";
    FD1P3AX intgOut3_i23 (.D(intgOut0_28__N_735[23]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i23.GSR = "ENABLED";
    FD1P3AX intgOut3_i24 (.D(intgOut0_28__N_735[24]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i24.GSR = "ENABLED";
    FD1P3AX intgOut3_i25 (.D(intgOut0_28__N_735[25]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i25.GSR = "ENABLED";
    FD1P3AX intgOut3_i26 (.D(intgOut0_28__N_735[26]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i26.GSR = "ENABLED";
    FD1P3AX intgOut3_i27 (.D(intgOut0_28__N_735[27]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i27.GSR = "ENABLED";
    FD1P3AX intgOut3_i28 (.D(intgOut0_28__N_735[28]), .SP(clk_N_683_enable_185), 
            .CK(clk_N_683), .Q(intgOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam intgOut3_i28.GSR = "ENABLED";
    FD1P3AX Out0_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i1.GSR = "ENABLED";
    FD1P3AX Out0_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i2.GSR = "ENABLED";
    FD1P3AX Out0_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i3.GSR = "ENABLED";
    FD1P3AX Out0_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i4.GSR = "ENABLED";
    FD1P3AX Out0_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i5.GSR = "ENABLED";
    FD1P3AX Out0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i6.GSR = "ENABLED";
    FD1P3AX Out0_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i7.GSR = "ENABLED";
    FD1P3AX Out0_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i8.GSR = "ENABLED";
    FD1P3AX Out0_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i9.GSR = "ENABLED";
    FD1P3AX Out0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i10.GSR = "ENABLED";
    FD1P3AX Out0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i11.GSR = "ENABLED";
    FD1P3AX Out0_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i12.GSR = "ENABLED";
    FD1P3AX Out0_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i13.GSR = "ENABLED";
    FD1P3AX Out0_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i14.GSR = "ENABLED";
    FD1P3AX Out0_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i15.GSR = "ENABLED";
    FD1P3AX Out0_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i16.GSR = "ENABLED";
    FD1P3AX Out0_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i17.GSR = "ENABLED";
    FD1P3AX Out0_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i18.GSR = "ENABLED";
    FD1P3AX Out0_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i19.GSR = "ENABLED";
    FD1P3AX Out0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i20.GSR = "ENABLED";
    FD1P3AX Out0_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i21.GSR = "ENABLED";
    FD1P3AX Out0_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i22.GSR = "ENABLED";
    FD1P3AX Out0_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i23.GSR = "ENABLED";
    FD1P3AX Out0_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i24.GSR = "ENABLED";
    FD1P3AX Out0_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i25.GSR = "ENABLED";
    FD1P3AX Out0_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i26.GSR = "ENABLED";
    FD1P3AX Out0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i27.GSR = "ENABLED";
    FD1P3AX Out0_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_213), 
            .CK(clk_N_683), .Q(Out0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out0_i28.GSR = "ENABLED";
    FD1P3AX Out1_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i1.GSR = "ENABLED";
    FD1P3AX Out1_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i2.GSR = "ENABLED";
    FD1P3AX Out1_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i3.GSR = "ENABLED";
    FD1P3AX Out1_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i4.GSR = "ENABLED";
    FD1P3AX Out1_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i5.GSR = "ENABLED";
    FD1P3AX Out1_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i6.GSR = "ENABLED";
    FD1P3AX Out1_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i7.GSR = "ENABLED";
    FD1P3AX Out1_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i8.GSR = "ENABLED";
    FD1P3AX Out1_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i9.GSR = "ENABLED";
    FD1P3AX Out1_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i10.GSR = "ENABLED";
    FD1P3AX Out1_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i11.GSR = "ENABLED";
    FD1P3AX Out1_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i12.GSR = "ENABLED";
    FD1P3AX Out1_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i13.GSR = "ENABLED";
    FD1P3AX Out1_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i14.GSR = "ENABLED";
    FD1P3AX Out1_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i15.GSR = "ENABLED";
    FD1P3AX Out1_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i16.GSR = "ENABLED";
    FD1P3AX Out1_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i17.GSR = "ENABLED";
    FD1P3AX Out1_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i18.GSR = "ENABLED";
    FD1P3AX Out1_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i19.GSR = "ENABLED";
    FD1P3AX Out1_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i20.GSR = "ENABLED";
    FD1P3AX Out1_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i21.GSR = "ENABLED";
    FD1P3AX Out1_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i22.GSR = "ENABLED";
    FD1P3AX Out1_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i23.GSR = "ENABLED";
    FD1P3AX Out1_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i24.GSR = "ENABLED";
    FD1P3AX Out1_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i25.GSR = "ENABLED";
    FD1P3AX Out1_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i26.GSR = "ENABLED";
    FD1P3AX Out1_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i27.GSR = "ENABLED";
    FD1P3AX Out1_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_241), 
            .CK(clk_N_683), .Q(Out1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out1_i28.GSR = "ENABLED";
    FD1P3AX Out2_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i1.GSR = "ENABLED";
    FD1P3AX Out2_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i2.GSR = "ENABLED";
    FD1P3AX Out2_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i3.GSR = "ENABLED";
    FD1P3AX Out2_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i4.GSR = "ENABLED";
    FD1P3AX Out2_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i5.GSR = "ENABLED";
    FD1P3AX Out2_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i6.GSR = "ENABLED";
    FD1P3AX Out2_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i7.GSR = "ENABLED";
    FD1P3AX Out2_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i8.GSR = "ENABLED";
    FD1P3AX Out2_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i9.GSR = "ENABLED";
    FD1P3AX Out2_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i10.GSR = "ENABLED";
    FD1P3AX Out2_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i11.GSR = "ENABLED";
    FD1P3AX Out2_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i12.GSR = "ENABLED";
    FD1P3AX Out2_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i13.GSR = "ENABLED";
    FD1P3AX Out2_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i14.GSR = "ENABLED";
    FD1P3AX Out2_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i15.GSR = "ENABLED";
    FD1P3AX Out2_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i16.GSR = "ENABLED";
    FD1P3AX Out2_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i17.GSR = "ENABLED";
    FD1P3AX Out2_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i18.GSR = "ENABLED";
    FD1P3AX Out2_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i19.GSR = "ENABLED";
    FD1P3AX Out2_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i20.GSR = "ENABLED";
    FD1P3AX Out2_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i21.GSR = "ENABLED";
    FD1P3AX Out2_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i22.GSR = "ENABLED";
    FD1P3AX Out2_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i23.GSR = "ENABLED";
    FD1P3AX Out2_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i24.GSR = "ENABLED";
    FD1P3AX Out2_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i25.GSR = "ENABLED";
    FD1P3AX Out2_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i26.GSR = "ENABLED";
    FD1P3AX Out2_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i27.GSR = "ENABLED";
    FD1P3AX Out2_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_269), 
            .CK(clk_N_683), .Q(Out2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out2_i28.GSR = "ENABLED";
    FD1P3AX Out3_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i1.GSR = "ENABLED";
    FD1P3AX Out3_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i2.GSR = "ENABLED";
    FD1P3AX Out3_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i3.GSR = "ENABLED";
    FD1P3AX Out3_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i4.GSR = "ENABLED";
    FD1P3AX Out3_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i5.GSR = "ENABLED";
    FD1P3AX Out3_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i6.GSR = "ENABLED";
    FD1P3AX Out3_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i7.GSR = "ENABLED";
    FD1P3AX Out3_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i8.GSR = "ENABLED";
    FD1P3AX Out3_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i9.GSR = "ENABLED";
    FD1P3AX Out3_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i10.GSR = "ENABLED";
    FD1P3AX Out3_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i11.GSR = "ENABLED";
    FD1P3AX Out3_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i12.GSR = "ENABLED";
    FD1P3AX Out3_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i13.GSR = "ENABLED";
    FD1P3AX Out3_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i14.GSR = "ENABLED";
    FD1P3AX Out3_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i15.GSR = "ENABLED";
    FD1P3AX Out3_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i16.GSR = "ENABLED";
    FD1P3AX Out3_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i17.GSR = "ENABLED";
    FD1P3AX Out3_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i18.GSR = "ENABLED";
    FD1P3AX Out3_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i19.GSR = "ENABLED";
    FD1P3AX Out3_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i20.GSR = "ENABLED";
    FD1P3AX Out3_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i21.GSR = "ENABLED";
    FD1P3AX Out3_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i22.GSR = "ENABLED";
    FD1P3AX Out3_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i23.GSR = "ENABLED";
    FD1P3AX Out3_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i24.GSR = "ENABLED";
    FD1P3AX Out3_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i25.GSR = "ENABLED";
    FD1P3AX Out3_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i26.GSR = "ENABLED";
    FD1P3AX Out3_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i27.GSR = "ENABLED";
    FD1P3AX Out3_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_297), 
            .CK(clk_N_683), .Q(Out3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam Out3_i28.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_325), 
            .CK(clk_N_683), .Q(backOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut2_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i1 (.D(backOut0_28__N_1416[1]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i2 (.D(backOut0_28__N_1416[2]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i3 (.D(backOut0_28__N_1416[3]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i4 (.D(backOut0_28__N_1416[4]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i5 (.D(backOut1_28__N_1445[5]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i6 (.D(backOut1_28__N_1445[6]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i7 (.D(backOut0_28__N_1416[7]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i8 (.D(backOut0_28__N_1416[8]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i9 (.D(backOut1_28__N_1445[9]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i10 (.D(backOut1_28__N_1445[10]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i11 (.D(backOut1_28__N_1445[11]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i12 (.D(backOut0_28__N_1416[12]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i13 (.D(backOut0_28__N_1416[13]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i14 (.D(backOut0_28__N_1416[14]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i15 (.D(backOut0_28__N_1416[15]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i16 (.D(backOut0_28__N_1416[16]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i17 (.D(backOut0_28__N_1416[17]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i18 (.D(backOut0_28__N_1416[18]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i19 (.D(backOut0_28__N_1416[19]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i20 (.D(backOut1_28__N_1445[20]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i21 (.D(backOut1_28__N_1445[21]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i22 (.D(backOut1_28__N_1445[22]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i23 (.D(backOut0_28__N_1416[23]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i24 (.D(backOut0_28__N_1416[24]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i25 (.D(backOut1_28__N_1445[25]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i26 (.D(backOut2_28__N_1474[26]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i27 (.D(backOut1_28__N_1445[27]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i28 (.D(backOut0_28__N_1416[28]), .SP(clk_N_683_enable_353), 
            .CK(clk_N_683), .Q(backOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam backOut3_i0_i28.GSR = "DISABLED";
    PFUMX mux_1193_i2 (.BLUT(n5091), .ALUT(n5049), .C0(n2436), .Z(n5139));
    LUT4 i1_2_lut_adj_57 (.A(Out0[8]), .B(Out0[12]), .Z(n6_adj_1832)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam i1_2_lut_adj_57.init = 16'heeee;
    PFUMX mux_1193_i1 (.BLUT(n5047), .ALUT(n5045), .C0(n2436), .Z(n5137));
    LUT4 i13930_4_lut_4_lut (.A(n920), .B(n3635), .C(addOut[19]), .D(n22208), 
         .Z(intgOut0_28__N_735[19])) /* synthesis lut_function=(!(A (D)+!A (B+((D)+!C)))) */ ;
    defparam i13930_4_lut_4_lut.init = 16'h00ba;
    LUT4 mux_1799_i15_4_lut (.A(\speed_m4[14] ), .B(\speed_m3[14] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i15_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut (.A(ss[3]), .B(n19740), .C(n22208), .D(n21565), .Z(clk_N_683_enable_41)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hc4c0;
    FD1S3AX subOut_i1 (.D(subOut_24__N_1135[1]), .CK(clk_N_683), .Q(subOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i1.GSR = "ENABLED";
    FD1S3AX subOut_i2 (.D(subOut_24__N_1135[2]), .CK(clk_N_683), .Q(subOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i2.GSR = "ENABLED";
    FD1S3AX subOut_i3 (.D(subOut_24__N_1135[3]), .CK(clk_N_683), .Q(subOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i3.GSR = "ENABLED";
    FD1S3AX subOut_i4 (.D(subOut_24__N_1135[4]), .CK(clk_N_683), .Q(subOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i4.GSR = "ENABLED";
    FD1S3AX subOut_i5 (.D(subOut_24__N_1135[5]), .CK(clk_N_683), .Q(subOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i5.GSR = "ENABLED";
    FD1S3AX subOut_i6 (.D(subOut_24__N_1135[6]), .CK(clk_N_683), .Q(subOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i6.GSR = "ENABLED";
    FD1S3AX subOut_i7 (.D(subOut_24__N_1135[7]), .CK(clk_N_683), .Q(subOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i7.GSR = "ENABLED";
    FD1S3AX subOut_i8 (.D(subOut_24__N_1135[8]), .CK(clk_N_683), .Q(subOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i8.GSR = "ENABLED";
    FD1S3AX subOut_i9 (.D(subOut_24__N_1135[9]), .CK(clk_N_683), .Q(subOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i9.GSR = "ENABLED";
    FD1S3AX subOut_i10 (.D(subOut_24__N_1135[10]), .CK(clk_N_683), .Q(subOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i10.GSR = "ENABLED";
    FD1S3AX subOut_i11 (.D(subOut_24__N_1135[11]), .CK(clk_N_683), .Q(subOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i11.GSR = "ENABLED";
    FD1S3AX subOut_i12 (.D(subOut_24__N_1135[12]), .CK(clk_N_683), .Q(subOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i12.GSR = "ENABLED";
    FD1S3AX subOut_i13 (.D(subOut_24__N_1135[13]), .CK(clk_N_683), .Q(subOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i13.GSR = "ENABLED";
    FD1S3AX subOut_i14 (.D(subOut_24__N_1135[14]), .CK(clk_N_683), .Q(subOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i14.GSR = "ENABLED";
    FD1S3AX subOut_i15 (.D(subOut_24__N_1135[15]), .CK(clk_N_683), .Q(subOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i15.GSR = "ENABLED";
    FD1S3AX subOut_i16 (.D(subOut_24__N_1135[16]), .CK(clk_N_683), .Q(subOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i16.GSR = "ENABLED";
    FD1S3AX subOut_i17 (.D(subOut_24__N_1135[17]), .CK(clk_N_683), .Q(subOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i17.GSR = "ENABLED";
    FD1S3AX subOut_i18 (.D(subOut_24__N_1135[18]), .CK(clk_N_683), .Q(subOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i18.GSR = "ENABLED";
    FD1S3AX subOut_i19 (.D(subOut_24__N_1135[19]), .CK(clk_N_683), .Q(subOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i19.GSR = "ENABLED";
    FD1S3AX subOut_i20 (.D(subOut_24__N_1135[20]), .CK(clk_N_683), .Q(subOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i20.GSR = "ENABLED";
    FD1S3AX subOut_i21 (.D(subOut_24__N_1135[21]), .CK(clk_N_683), .Q(subOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i21.GSR = "ENABLED";
    FD1S3AX subOut_i23 (.D(subOut_24__N_1135[24]), .CK(clk_N_683), .Q(subOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam subOut_i23.GSR = "ENABLED";
    LUT4 mux_205_i4_3_lut_4_lut_3_lut (.A(n30_adj_1833), .B(n1166[15]), 
         .C(n2164[3]), .Z(n1302[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(334[25:42])
    defparam mux_205_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_205_i8_3_lut_4_lut_3_lut (.A(n30_adj_1833), .B(n1166[15]), 
         .C(n2164[7]), .Z(n1302[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(334[25:42])
    defparam mux_205_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_205_i10_3_lut_4_lut_3_lut (.A(n30_adj_1833), .B(n1166[15]), 
         .C(n2164[9]), .Z(n1302[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(334[25:42])
    defparam mux_205_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 n9_bdd_4_lut (.A(n21528), .B(n21550), .C(ss[0]), .D(ss[1]), 
         .Z(n15941)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))) */ ;
    defparam n9_bdd_4_lut.init = 16'ha88a;
    LUT4 mux_205_i9_3_lut_4_lut_3_lut (.A(n30_adj_1833), .B(n1166[15]), 
         .C(n2164[8]), .Z(n1302[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(334[25:42])
    defparam mux_205_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 ss_1__bdd_4_lut_18293 (.A(n22208), .B(ss[0]), .C(ss[2]), .D(ss[3]), 
         .Z(n16618)) /* synthesis lut_function=(A+(B+(C (D)+!C !(D)))) */ ;
    defparam ss_1__bdd_4_lut_18293.init = 16'hfeef;
    LUT4 mux_1799_i14_4_lut (.A(\speed_m4[13] ), .B(\speed_m3[13] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i14_4_lut.init = 16'hcac0;
    LUT4 mux_205_i7_3_lut_4_lut_3_lut (.A(n30_adj_1833), .B(n1166[15]), 
         .C(n2164[6]), .Z(n1302[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(334[25:42])
    defparam mux_205_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_205_i6_3_lut_4_lut_3_lut (.A(n30_adj_1833), .B(n1166[15]), 
         .C(n2164[5]), .Z(n1302[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(334[25:42])
    defparam mux_205_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_212_i4_3_lut_4_lut_3_lut (.A(n30), .B(n1187[15]), .C(n2176[3]), 
         .Z(n1346[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(342[25:42])
    defparam mux_212_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_1799_i12_4_lut (.A(\speed_m4[11] ), .B(\speed_m3[11] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i12_4_lut.init = 16'hcac0;
    LUT4 mux_212_i8_3_lut_4_lut_3_lut (.A(n30), .B(n1187[15]), .C(n2176[7]), 
         .Z(n1346[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(342[25:42])
    defparam mux_212_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i5_4_lut (.A(n9), .B(n7_c), .C(n1208[10]), .D(n1208[13]), .Z(n30_adj_1834)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i3_2_lut (.A(n1208[14]), .B(n1208[12]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_58 (.A(n1208[11]), .B(n1208[9]), .C(n10_adj_1835), 
         .D(n1208[7]), .Z(n7_c)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_58.init = 16'haaa8;
    LUT4 mux_212_i10_3_lut_4_lut_3_lut (.A(n30), .B(n1187[15]), .C(n2176[9]), 
         .Z(n1346[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(342[25:42])
    defparam mux_212_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i4_4_lut_adj_59 (.A(n1208[6]), .B(n8), .C(n1208[4]), .D(n4), 
         .Z(n10_adj_1835)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_59.init = 16'hfeee;
    LUT4 mux_212_i9_3_lut_4_lut_3_lut (.A(n30), .B(n1187[15]), .C(n2176[8]), 
         .Z(n1346[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(342[25:42])
    defparam mux_212_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_212_i7_3_lut_4_lut_3_lut (.A(n30), .B(n1187[15]), .C(n2176[6]), 
         .Z(n1346[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(342[25:42])
    defparam mux_212_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i2_2_lut_adj_60 (.A(n1208[5]), .B(n1208[8]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_60.init = 16'heeee;
    LUT4 i1_4_lut_adj_61 (.A(n1208[3]), .B(n1208[2]), .C(n1208[1]), .D(n1208[0]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_61.init = 16'haaa8;
    PFUMX i3392 (.BLUT(n2484[1]), .ALUT(n5688), .C0(n21483), .Z(n5689));
    LUT4 mux_212_i6_3_lut_4_lut_3_lut (.A(n30), .B(n1187[15]), .C(n2176[5]), 
         .Z(n1346[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(342[25:42])
    defparam mux_212_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i10236_3_lut_4_lut (.A(n1208[15]), .B(n30_adj_1834), .C(n18815), 
         .D(clk_N_683_enable_392), .Z(n12666)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(350[7:42])
    defparam i10236_3_lut_4_lut.init = 16'hf700;
    LUT4 mux_1799_i11_4_lut (.A(\speed_m4[10] ), .B(\speed_m3[10] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i11_4_lut.init = 16'hcac0;
    PFUMX i3394 (.BLUT(n2484[2]), .ALUT(n5690), .C0(n21483), .Z(n5691));
    LUT4 mux_1799_i7_4_lut (.A(\speed_m4[6] ), .B(\speed_m3[6] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i7_4_lut.init = 16'hcac0;
    LUT4 mux_219_i4_3_lut_4_lut_3_lut (.A(n30_adj_1834), .B(n1208[15]), 
         .C(n2188[3]), .Z(n1390[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(350[25:42])
    defparam mux_219_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i14184_2_lut_rep_279_4_lut (.A(n21526), .B(n21577), .C(n21578), 
         .D(n56), .Z(n21488)) /* synthesis lut_function=(A (B+(C+(D)))+!A (D)) */ ;
    defparam i14184_2_lut_rep_279_4_lut.init = 16'hffa8;
    LUT4 i59_2_lut_4_lut (.A(n21526), .B(n21577), .C(n21578), .D(n56), 
         .Z(n57)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(D))) */ ;
    defparam i59_2_lut_4_lut.init = 16'h5700;
    LUT4 i1_2_lut_rep_374 (.A(ss[0]), .B(ss[2]), .Z(n21583)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_374.init = 16'h8888;
    LUT4 mux_219_i10_3_lut_4_lut_3_lut (.A(n30_adj_1834), .B(n1208[15]), 
         .C(n2188[9]), .Z(n1390[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(350[25:42])
    defparam mux_219_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i1_2_lut_rep_356_3_lut (.A(ss[0]), .B(ss[2]), .C(ss[1]), .Z(n21565)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_356_3_lut.init = 16'h8080;
    LUT4 i8797_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[2]), .C(ss[3]), .D(ss[1]), 
         .Z(n15)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i8797_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i13686_2_lut_rep_375 (.A(ss[0]), .B(ss[1]), .Z(n21584)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13686_2_lut_rep_375.init = 16'h8888;
    LUT4 i7789_2_lut_3_lut (.A(ss[0]), .B(ss[1]), .C(ss[2]), .Z(n14)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i7789_2_lut_3_lut.init = 16'h7878;
    LUT4 mux_1799_i6_4_lut (.A(\speed_m4[5] ), .B(\speed_m3[5] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i6_4_lut.init = 16'hcac0;
    CCU2D sub_16_rep_3_add_2_9 (.A0(subIn2[7]), .B0(n16648), .C0(n16541), 
          .D0(n5701), .A1(subIn2[8]), .B1(n16648), .C1(n16541), .D1(n5703), 
          .CIN(n18638), .COUT(n18639), .S0(n27[7]), .S1(n27[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_9.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_9.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(n21569), .B(n22208), .C(n21565), .D(ss[3]), 
         .Z(clk_N_683_enable_297)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam i1_4_lut_4_lut.init = 16'hb888;
    CCU2D add_15798_4 (.A0(addOut[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18707), .COUT(n18708));
    defparam add_15798_4.INIT0 = 16'h5aaa;
    defparam add_15798_4.INIT1 = 16'h5555;
    defparam add_15798_4.INJECT1_0 = "NO";
    defparam add_15798_4.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_adj_62 (.A(n21569), .B(n22208), .C(n19776), .D(ss[1]), 
         .Z(clk_N_683_enable_185)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(B+(C+!(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_62.init = 16'h8b88;
    LUT4 mux_1799_i5_4_lut (.A(\speed_m4[4] ), .B(\speed_m3[4] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i5_4_lut.init = 16'hcac0;
    PFUMX i3396 (.BLUT(n2484[3]), .ALUT(n5692), .C0(n21483), .Z(n5693));
    LUT4 i1_4_lut_4_lut_adj_63 (.A(n21569), .B(n22208), .C(n19776), .D(ss[1]), 
         .Z(clk_N_683_enable_157)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+(C+(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_63.init = 16'h888b;
    LUT4 mux_219_i7_3_lut_4_lut_3_lut (.A(n30_adj_1834), .B(n1208[15]), 
         .C(n2188[6]), .Z(n1390[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(350[25:42])
    defparam mux_219_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i1_4_lut_4_lut_adj_64 (.A(n21569), .B(n22208), .C(n19779), .D(n21601), 
         .Z(clk_N_683_enable_213)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+(C+(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_64.init = 16'h888b;
    LUT4 mux_1799_i3_4_lut (.A(\speed_m4[2] ), .B(\speed_m3[2] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i3_4_lut.init = 16'hcac0;
    PFUMX i3398 (.BLUT(n2484[4]), .ALUT(n5694), .C0(n21483), .Z(n5695));
    LUT4 i1_4_lut_4_lut_adj_65 (.A(n21569), .B(n22208), .C(n19897), .D(n21601), 
         .Z(clk_N_683_enable_269)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B+((D)+!C))) */ ;
    defparam i1_4_lut_4_lut_adj_65.init = 16'h88b8;
    LUT4 i3433_2_lut_rep_377 (.A(n22208), .B(n22203), .Z(clk_N_683_enable_392)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam i3433_2_lut_rep_377.init = 16'h8888;
    LUT4 mux_1799_i2_4_lut (.A(\speed_m4[1] ), .B(\speed_m3[1] ), .C(n21544), 
         .D(n4132), .Z(subIn2_24__N_1301[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(147[18] 151[17])
    defparam mux_1799_i2_4_lut.init = 16'hcac0;
    LUT4 i17974_2_lut_3_lut_4_lut_4_lut (.A(n21548), .B(n21508), .C(n21549), 
         .D(n21552), .Z(multIn2[4])) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i17974_2_lut_3_lut_4_lut_4_lut.init = 16'h1115;
    CCU2D sub_16_rep_3_add_2_7 (.A0(subIn2[5]), .B0(n16648), .C0(n16541), 
          .D0(n5697), .A1(subIn2[6]), .B1(n16648), .C1(n16541), .D1(n5699), 
          .CIN(n18637), .COUT(n18638), .S0(n27[5]), .S1(n27[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_7.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_7.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_5 (.A0(subIn2[3]), .B0(n16648), .C0(n16541), 
          .D0(n5693), .A1(subIn2[4]), .B1(n16648), .C1(n16541), .D1(n5695), 
          .CIN(n18636), .COUT(n18637), .S0(n27[3]), .S1(n27[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_5.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_5.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_5.INJECT1_1 = "NO";
    CCU2D add_15798_2 (.A0(addOut[7]), .B0(addOut[6]), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18707));
    defparam add_15798_2.INIT0 = 16'h1000;
    defparam add_15798_2.INIT1 = 16'h5555;
    defparam add_15798_2.INJECT1_0 = "NO";
    defparam add_15798_2.INJECT1_1 = "NO";
    PFUMX i3400 (.BLUT(n2484[5]), .ALUT(n5696), .C0(n21483), .Z(n5697));
    LUT4 i1_4_lut_4_lut_else_4_lut (.A(ss[1]), .B(ss[2]), .C(ss[3]), .D(ss[0]), 
         .Z(n21609)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_else_4_lut.init = 16'h4000;
    LUT4 i2_3_lut_rep_299_4_lut (.A(n21577), .B(n21549), .C(n21529), .D(n21528), 
         .Z(n21508)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(174[9:17])
    defparam i2_3_lut_rep_299_4_lut.init = 16'he000;
    LUT4 mux_136_i1_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[0]), 
         .D(backOut1[0]), .Z(n588[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i25_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[24]), 
         .D(backOut1[24]), .Z(n588[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i27_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[26]), 
         .D(backOut1[26]), .Z(n588[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10366_2_lut_3_lut_4_lut (.A(n22208), .B(n22203), .C(n21607), 
         .D(n21608), .Z(n12641)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam i10366_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 mux_136_i28_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[27]), 
         .D(backOut1[27]), .Z(n588[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i28_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3402 (.BLUT(n2484[6]), .ALUT(n5698), .C0(n21483), .Z(n5699));
    LUT4 mux_136_i26_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[25]), 
         .D(backOut1[25]), .Z(n588[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i26_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3404 (.BLUT(n2484[7]), .ALUT(n5700), .C0(n21483), .Z(n5701));
    LUT4 mux_136_i24_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[23]), 
         .D(backOut1[23]), .Z(n588[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i18_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[17]), 
         .D(backOut1[17]), .Z(n588[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i23_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[22]), 
         .D(backOut1[22]), .Z(n588[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i23_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3406 (.BLUT(n2484[8]), .ALUT(n5702), .C0(n21483), .Z(n5703));
    LUT4 mux_136_i29_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[28]), 
         .D(backOut1[28]), .Z(n588[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i29_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3408 (.BLUT(n2484[9]), .ALUT(n5704), .C0(n21483), .Z(n5705));
    LUT4 mux_136_i22_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[21]), 
         .D(backOut1[21]), .Z(n588[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i22_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3410 (.BLUT(n2484[10]), .ALUT(n5706), .C0(n21483), .Z(n5707));
    PFUMX i3412 (.BLUT(n2484[11]), .ALUT(n5708), .C0(n21483), .Z(n5709));
    LUT4 mux_136_i21_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[20]), 
         .D(backOut1[20]), .Z(n588[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i20_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[19]), 
         .D(backOut1[19]), .Z(n588[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i19_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[18]), 
         .D(backOut1[18]), .Z(n588[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i19_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3414 (.BLUT(n2484[12]), .ALUT(n5710), .C0(n21483), .Z(n5711));
    LUT4 mux_136_i9_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[8]), 
         .D(backOut1[8]), .Z(n588[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i2_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[1]), 
         .D(backOut1[1]), .Z(n588[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i2_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3416 (.BLUT(n2484[13]), .ALUT(n5712), .C0(n21483), .Z(n5713));
    CCU2D add_15799_29 (.A0(addOut[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18706), 
          .S1(n3635));
    defparam add_15799_29.INIT0 = 16'h5aaa;
    defparam add_15799_29.INIT1 = 16'h0000;
    defparam add_15799_29.INJECT1_0 = "NO";
    defparam add_15799_29.INJECT1_1 = "NO";
    LUT4 mux_136_i10_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[9]), 
         .D(backOut1[9]), .Z(n588[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i17_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[16]), 
         .D(backOut1[16]), .Z(n588[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i17_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3418 (.BLUT(n2484[14]), .ALUT(n5714), .C0(n21483), .Z(n5715));
    LUT4 mux_136_i3_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[2]), 
         .D(backOut1[2]), .Z(n588[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i3_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15799_27 (.A0(addOut[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18705), .COUT(n18706));
    defparam add_15799_27.INIT0 = 16'h0aaa;
    defparam add_15799_27.INIT1 = 16'h0aaa;
    defparam add_15799_27.INJECT1_0 = "NO";
    defparam add_15799_27.INJECT1_1 = "NO";
    LUT4 mux_136_i7_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[6]), 
         .D(backOut1[6]), .Z(n588[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i12_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[11]), 
         .D(backOut1[11]), .Z(n588[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i11_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[10]), 
         .D(backOut1[10]), .Z(n588[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i8_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[7]), 
         .D(backOut1[7]), .Z(n588[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i8_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3420 (.BLUT(n2484[15]), .ALUT(n5716), .C0(n21483), .Z(n5717));
    LUT4 mux_136_i13_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[12]), 
         .D(backOut1[12]), .Z(n588[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i5_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[4]), 
         .D(backOut1[4]), .Z(n588[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i5_3_lut_4_lut.init = 16'hfd20;
    PFUMX i3422 (.BLUT(n2484[16]), .ALUT(n5718), .C0(n21483), .Z(n5719));
    LUT4 mux_136_i4_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[3]), 
         .D(backOut1[3]), .Z(n588[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_219_i9_3_lut_4_lut_3_lut (.A(n30_adj_1834), .B(n1208[15]), 
         .C(n2188[8]), .Z(n1390[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(350[25:42])
    defparam mux_219_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    PFUMX i3424 (.BLUT(n2484[17]), .ALUT(n5720), .C0(n21483), .Z(n5721));
    LUT4 mux_136_i15_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[14]), 
         .D(backOut1[14]), .Z(n588[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i14_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[13]), 
         .D(backOut1[13]), .Z(n588[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_219_i8_3_lut_4_lut_3_lut (.A(n30_adj_1834), .B(n1208[15]), 
         .C(n2188[7]), .Z(n1390[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(350[25:42])
    defparam mux_219_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_136_i6_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[5]), 
         .D(backOut1[5]), .Z(n588[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i16_3_lut_4_lut (.A(n21584), .B(n21554), .C(backOut0[15]), 
         .D(backOut1[15]), .Z(n588[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(173[9:17])
    defparam mux_136_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_290_4_lut_4_lut (.A(n21551), .B(n21550), .C(n21577), 
         .D(n21529), .Z(n21499)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_290_4_lut_4_lut.init = 16'h5400;
    LUT4 mux_219_i6_3_lut_4_lut_3_lut (.A(n30_adj_1834), .B(n1208[15]), 
         .C(n2188[5]), .Z(n1390[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(350[25:42])
    defparam mux_219_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i14360_2_lut_rep_280_3_lut_3_lut (.A(n21551), .B(n42), .C(n21509), 
         .Z(n21489)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(165[9:16])
    defparam i14360_2_lut_rep_280_3_lut_3_lut.init = 16'hdcdc;
    PFUMX i3426 (.BLUT(n2484[18]), .ALUT(n5722), .C0(n21483), .Z(n5723));
    LUT4 i1_2_lut_rep_281_3_lut_3_lut (.A(n21551), .B(n42), .C(n21509), 
         .Z(n21490)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_281_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_3_lut_4_lut (.A(n22208), .B(n920), .C(addOut[7]), .D(n3635), 
         .Z(intgOut0_28__N_735[7])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1110;
    LUT4 i3_4_lut_4_lut (.A(n21485), .B(n21488), .C(n21500), .D(n21489), 
         .Z(n16648)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut_4_lut.init = 16'h0400;
    LUT4 i1_3_lut_4_lut_adj_66 (.A(n22208), .B(n920), .C(addOut[8]), .D(n3635), 
         .Z(intgOut0_28__N_735[8])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_66.init = 16'h1110;
    LUT4 i1_3_lut_4_lut_adj_67 (.A(n22208), .B(n920), .C(addOut[10]), 
         .D(n3635), .Z(intgOut0_28__N_735[10])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_67.init = 16'h1110;
    LUT4 i1_3_lut_4_lut_adj_68 (.A(n22208), .B(n920), .C(addOut[11]), 
         .D(n3635), .Z(intgOut0_28__N_735[11])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_68.init = 16'h1110;
    LUT4 mux_1800_i1_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[0] ), 
         .D(\speed_m2[0] ), .Z(subIn2_24__N_1114[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut_adj_69 (.A(n22208), .B(n920), .C(addOut[12]), 
         .D(n3635), .Z(intgOut0_28__N_735[12])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_69.init = 16'h1110;
    LUT4 mux_1800_i19_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[18] ), 
         .D(\speed_m2[18] ), .Z(subIn2_24__N_1114[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i18_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[17] ), 
         .D(\speed_m2[17] ), .Z(subIn2_24__N_1114[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i17_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[16] ), 
         .D(\speed_m2[16] ), .Z(subIn2_24__N_1114[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i16_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[15] ), 
         .D(\speed_m2[15] ), .Z(subIn2_24__N_1114[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i15_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[14] ), 
         .D(\speed_m2[14] ), .Z(subIn2_24__N_1114[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i15_3_lut_4_lut.init = 16'hfb40;
    PFUMX i3428 (.BLUT(n2484[19]), .ALUT(n5724), .C0(n21483), .Z(n5725));
    CCU2D add_191_11 (.A0(Out3[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18443), 
          .COUT(n18444), .S0(n1208[9]), .S1(n1208[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_11.INIT0 = 16'h5aaa;
    defparam add_191_11.INIT1 = 16'h5aaa;
    defparam add_191_11.INJECT1_0 = "NO";
    defparam add_191_11.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_3 (.A0(subIn2[1]), .B0(n16648), .C0(n16541), 
          .D0(n5689), .A1(subIn2[2]), .B1(n16648), .C1(n16541), .D1(n5691), 
          .CIN(n18635), .COUT(n18636), .S0(n27[1]), .S1(n27[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_3.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_3.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_3.INJECT1_1 = "NO";
    LUT4 mux_1800_i14_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[13] ), 
         .D(\speed_m2[13] ), .Z(subIn2_24__N_1114[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i14_3_lut_4_lut.init = 16'hfb40;
    CCU2D sub_16_rep_3_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(subIn2[0]), .B1(n16648), .C1(n16541), .D1(n5254), 
          .COUT(n18635), .S1(n27[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_1.INIT0 = 16'h0000;
    defparam sub_16_rep_3_add_2_1.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_1.INJECT1_1 = "NO";
    CCU2D add_15799_25 (.A0(addOut[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18704), .COUT(n18705));
    defparam add_15799_25.INIT0 = 16'h0aaa;
    defparam add_15799_25.INIT1 = 16'h0aaa;
    defparam add_15799_25.INJECT1_0 = "NO";
    defparam add_15799_25.INJECT1_1 = "NO";
    LUT4 mux_1800_i12_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[11] ), 
         .D(\speed_m2[11] ), .Z(subIn2_24__N_1114[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i12_3_lut_4_lut.init = 16'hfb40;
    PFUMX i3432 (.BLUT(n2484[20]), .ALUT(n5728), .C0(n21483), .Z(n5729));
    LUT4 i1_3_lut_4_lut_adj_70 (.A(n22208), .B(n920), .C(addOut[13]), 
         .D(n3635), .Z(intgOut0_28__N_735[13])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_70.init = 16'h1110;
    PFUMX i2960 (.BLUT(n2484[0]), .ALUT(n5253), .C0(n21483), .Z(n5254));
    LUT4 mux_1800_i11_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[10] ), 
         .D(\speed_m2[10] ), .Z(subIn2_24__N_1114[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i7_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[6] ), 
         .D(\speed_m2[6] ), .Z(subIn2_24__N_1114[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i6_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[5] ), 
         .D(\speed_m2[5] ), .Z(subIn2_24__N_1114[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1800_i5_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[4] ), 
         .D(\speed_m2[4] ), .Z(subIn2_24__N_1114[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i5_3_lut_4_lut.init = 16'hfb40;
    PFUMX addIn2_28__I_29_i29 (.BLUT(n618[28]), .ALUT(addIn2_28__N_1337[28]), 
          .C0(n20447), .Z(addIn2_28__N_1207[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D addOut_2063_add_4_29 (.A0(multOut[27]), .B0(n16618), .C0(addOut[27]), 
          .D0(addIn2_28__N_1207[27]), .A1(multOut[28]), .B1(n16618), .C1(addOut[28]), 
          .D1(addIn2_28__N_1207[28]), .CIN(n18570), .S0(n121[27]), .S1(n121[28]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_29.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_29.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_29.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_29.INJECT1_1 = "NO";
    CCU2D add_191_9 (.A0(Out3[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18442), 
          .COUT(n18443), .S0(n1208[7]), .S1(n1208[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_9.INIT0 = 16'h5aaa;
    defparam add_191_9.INIT1 = 16'h5aaa;
    defparam add_191_9.INJECT1_0 = "NO";
    defparam add_191_9.INJECT1_1 = "NO";
    LUT4 mux_1800_i3_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[2] ), 
         .D(\speed_m2[2] ), .Z(subIn2_24__N_1114[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i3_3_lut_4_lut.init = 16'hfb40;
    PFUMX addIn2_28__I_29_i28 (.BLUT(n618[27]), .ALUT(addIn2_28__N_1337[27]), 
          .C0(n20447), .Z(addIn2_28__N_1207[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1179_17 (.A0(n5167), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5169), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18411), 
          .COUT(n18412), .S0(n2244[15]), .S1(n2244[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_17.INIT0 = 16'hf555;
    defparam add_1179_17.INIT1 = 16'hf555;
    defparam add_1179_17.INJECT1_0 = "NO";
    defparam add_1179_17.INJECT1_1 = "NO";
    CCU2D add_1179_15 (.A0(n5163), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5165), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18410), 
          .COUT(n18411), .S0(n2244[13]), .S1(n2244[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_15.INIT0 = 16'hf555;
    defparam add_1179_15.INIT1 = 16'hf555;
    defparam add_1179_15.INJECT1_0 = "NO";
    defparam add_1179_15.INJECT1_1 = "NO";
    CCU2D add_1179_13 (.A0(n5159), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5161), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18409), 
          .COUT(n18410), .S0(n2244[11]), .S1(n2244[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_13.INIT0 = 16'hf555;
    defparam add_1179_13.INIT1 = 16'hf555;
    defparam add_1179_13.INJECT1_0 = "NO";
    defparam add_1179_13.INJECT1_1 = "NO";
    CCU2D add_1179_11 (.A0(n5155), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5157), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18408), 
          .COUT(n18409), .S0(n2244[9]), .S1(n2244[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_11.INIT0 = 16'hf555;
    defparam add_1179_11.INIT1 = 16'hf555;
    defparam add_1179_11.INJECT1_0 = "NO";
    defparam add_1179_11.INJECT1_1 = "NO";
    CCU2D add_1179_9 (.A0(n5151), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5153), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18407), 
          .COUT(n18408), .S0(n2244[7]), .S1(n2244[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_9.INIT0 = 16'hf555;
    defparam add_1179_9.INIT1 = 16'hf555;
    defparam add_1179_9.INJECT1_0 = "NO";
    defparam add_1179_9.INJECT1_1 = "NO";
    CCU2D add_1179_7 (.A0(n5147), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5149), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18406), 
          .COUT(n18407), .S0(n2244[5]), .S1(n2244[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_7.INIT0 = 16'hf555;
    defparam add_1179_7.INIT1 = 16'hf555;
    defparam add_1179_7.INJECT1_0 = "NO";
    defparam add_1179_7.INJECT1_1 = "NO";
    CCU2D add_1179_5 (.A0(n5143), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5145), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18405), 
          .COUT(n18406), .S0(n2244[3]), .S1(n2244[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_5.INIT0 = 16'hf555;
    defparam add_1179_5.INIT1 = 16'hf555;
    defparam add_1179_5.INJECT1_0 = "NO";
    defparam add_1179_5.INJECT1_1 = "NO";
    CCU2D add_1179_3 (.A0(n5139), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5141), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18404), 
          .COUT(n18405), .S0(n2244[1]), .S1(n2244[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_3.INIT0 = 16'hf555;
    defparam add_1179_3.INIT1 = 16'hf555;
    defparam add_1179_3.INJECT1_0 = "NO";
    defparam add_1179_3.INJECT1_1 = "NO";
    CCU2D add_1173_5 (.A0(n1145[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18400), 
          .COUT(n18401), .S0(n2152[3]), .S1(n2152[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(327[20:29])
    defparam add_1173_5.INIT0 = 16'hf555;
    defparam add_1173_5.INIT1 = 16'hf555;
    defparam add_1173_5.INJECT1_0 = "NO";
    defparam add_1173_5.INJECT1_1 = "NO";
    CCU2D add_1173_9 (.A0(n1145[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18402), 
          .COUT(n18403), .S0(n2152[7]), .S1(n2152[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(327[20:29])
    defparam add_1173_9.INIT0 = 16'hf555;
    defparam add_1173_9.INIT1 = 16'hf555;
    defparam add_1173_9.INJECT1_0 = "NO";
    defparam add_1173_9.INJECT1_1 = "NO";
    CCU2D add_1173_3 (.A0(n1145[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18399), 
          .COUT(n18400), .S0(n2152[1]), .S1(n2152[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(327[20:29])
    defparam add_1173_3.INIT0 = 16'hf555;
    defparam add_1173_3.INIT1 = 16'hf555;
    defparam add_1173_3.INJECT1_0 = "NO";
    defparam add_1173_3.INJECT1_1 = "NO";
    CCU2D add_1179_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5137), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18404), 
          .S1(n2244[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_1.INIT0 = 16'hF000;
    defparam add_1179_1.INIT1 = 16'h0aaa;
    defparam add_1179_1.INJECT1_0 = "NO";
    defparam add_1179_1.INJECT1_1 = "NO";
    CCU2D add_1173_7 (.A0(n1145[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18401), 
          .COUT(n18402), .S0(n2152[5]), .S1(n2152[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(327[20:29])
    defparam add_1173_7.INIT0 = 16'hf555;
    defparam add_1173_7.INIT1 = 16'hf555;
    defparam add_1173_7.INJECT1_0 = "NO";
    defparam add_1173_7.INJECT1_1 = "NO";
    CCU2D add_1173_11 (.A0(n1145[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18403), 
          .S0(n2152[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(327[20:29])
    defparam add_1173_11.INIT0 = 16'hf555;
    defparam add_1173_11.INIT1 = 16'h0000;
    defparam add_1173_11.INJECT1_0 = "NO";
    defparam add_1173_11.INJECT1_1 = "NO";
    CCU2D add_1173_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1145[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18399), 
          .S1(n2152[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(327[20:29])
    defparam add_1173_1.INIT0 = 16'hF000;
    defparam add_1173_1.INIT1 = 16'h0aaa;
    defparam add_1173_1.INJECT1_0 = "NO";
    defparam add_1173_1.INJECT1_1 = "NO";
    LUT4 mux_1800_i2_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[1] ), 
         .D(\speed_m2[1] ), .Z(subIn2_24__N_1114[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i2_3_lut_4_lut.init = 16'hfb40;
    CCU2D addOut_2063_add_4_27 (.A0(multOut[25]), .B0(n16618), .C0(addOut[25]), 
          .D0(addIn2_28__N_1207[25]), .A1(multOut[26]), .B1(n16618), .C1(addOut[26]), 
          .D1(addIn2_28__N_1207[26]), .CIN(n18569), .COUT(n18570), .S0(n121[25]), 
          .S1(n121[26]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_27.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_27.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_27.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_27.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_25 (.A0(multOut[23]), .B0(n16618), .C0(addOut[23]), 
          .D0(addIn2_28__N_1207[23]), .A1(multOut[24]), .B1(n16618), .C1(addOut[24]), 
          .D1(addIn2_28__N_1207[24]), .CIN(n18568), .COUT(n18569), .S0(n121[23]), 
          .S1(n121[24]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_25.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_25.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_25.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_25.INJECT1_1 = "NO";
    CCU2D add_15799_23 (.A0(addOut[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18703), .COUT(n18704));
    defparam add_15799_23.INIT0 = 16'h0aaa;
    defparam add_15799_23.INIT1 = 16'h0aaa;
    defparam add_15799_23.INJECT1_0 = "NO";
    defparam add_15799_23.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_23 (.A0(multOut[21]), .B0(n16618), .C0(addOut[21]), 
          .D0(addIn2_28__N_1207[21]), .A1(multOut[22]), .B1(n16618), .C1(addOut[22]), 
          .D1(addIn2_28__N_1207[22]), .CIN(n18567), .COUT(n18568), .S0(n121[21]), 
          .S1(n121[22]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_23.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_23.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_23.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_23.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_21 (.A0(multOut[19]), .B0(n16618), .C0(addOut[19]), 
          .D0(addIn2_28__N_1207[19]), .A1(multOut[20]), .B1(n16618), .C1(addOut[20]), 
          .D1(addIn2_28__N_1207[20]), .CIN(n18566), .COUT(n18567), .S0(n121[19]), 
          .S1(n121[20]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_21.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_21.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_21.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_21.INJECT1_1 = "NO";
    LUT4 i13582_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[19] ), 
         .D(\speed_m2[19] ), .Z(n5)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13582_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_15799_21 (.A0(addOut[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18702), .COUT(n18703));
    defparam add_15799_21.INIT0 = 16'h0aaa;
    defparam add_15799_21.INIT1 = 16'h0aaa;
    defparam add_15799_21.INJECT1_0 = "NO";
    defparam add_15799_21.INJECT1_1 = "NO";
    LUT4 mux_1800_i13_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[12] ), 
         .D(subIn2_24__N_1301[12]), .Z(subIn2_24__N_1114[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i13_3_lut_4_lut.init = 16'hfb40;
    PFUMX addIn2_28__I_29_i27 (.BLUT(n618[26]), .ALUT(addIn2_28__N_1337[26]), 
          .C0(n20447), .Z(addIn2_28__N_1207[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_1800_i10_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[9] ), 
         .D(subIn2_24__N_1301[9]), .Z(subIn2_24__N_1114[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i10_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_191_7 (.A0(Out3[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18441), 
          .COUT(n18442), .S0(n1208[5]), .S1(n1208[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_7.INIT0 = 16'h5aaa;
    defparam add_191_7.INIT1 = 16'h5aaa;
    defparam add_191_7.INJECT1_0 = "NO";
    defparam add_191_7.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i26 (.BLUT(n618[25]), .ALUT(addIn2_28__N_1337[25]), 
          .C0(n20447), .Z(addIn2_28__N_1207[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_1800_i9_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[8] ), 
         .D(subIn2_24__N_1301[8]), .Z(subIn2_24__N_1114[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i9_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_15799_19 (.A0(addOut[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18701), .COUT(n18702));
    defparam add_15799_19.INIT0 = 16'hf555;
    defparam add_15799_19.INIT1 = 16'hf555;
    defparam add_15799_19.INJECT1_0 = "NO";
    defparam add_15799_19.INJECT1_1 = "NO";
    CCU2D add_15799_17 (.A0(addOut[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18700), .COUT(n18701));
    defparam add_15799_17.INIT0 = 16'hf555;
    defparam add_15799_17.INIT1 = 16'hf555;
    defparam add_15799_17.INJECT1_0 = "NO";
    defparam add_15799_17.INJECT1_1 = "NO";
    CCU2D add_1176_11 (.A0(n1208[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18516), 
          .S0(n2188[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(351[20:29])
    defparam add_1176_11.INIT0 = 16'hf555;
    defparam add_1176_11.INIT1 = 16'h0000;
    defparam add_1176_11.INJECT1_0 = "NO";
    defparam add_1176_11.INJECT1_1 = "NO";
    CCU2D add_1176_9 (.A0(n1208[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18515), 
          .COUT(n18516), .S0(n2188[7]), .S1(n2188[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(351[20:29])
    defparam add_1176_9.INIT0 = 16'hf555;
    defparam add_1176_9.INIT1 = 16'hf555;
    defparam add_1176_9.INJECT1_0 = "NO";
    defparam add_1176_9.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i25 (.BLUT(n618[24]), .ALUT(addIn2_28__N_1337[24]), 
          .C0(n20447), .Z(addIn2_28__N_1207[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_1800_i8_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[7] ), 
         .D(subIn2_24__N_1301[7]), .Z(subIn2_24__N_1114[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i8_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_1176_7 (.A0(n1208[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18514), 
          .COUT(n18515), .S0(n2188[5]), .S1(n2188[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(351[20:29])
    defparam add_1176_7.INIT0 = 16'hf555;
    defparam add_1176_7.INIT1 = 16'hf555;
    defparam add_1176_7.INJECT1_0 = "NO";
    defparam add_1176_7.INJECT1_1 = "NO";
    CCU2D add_1176_5 (.A0(n1208[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18513), 
          .COUT(n18514), .S0(n2188[3]), .S1(n2188[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(351[20:29])
    defparam add_1176_5.INIT0 = 16'hf555;
    defparam add_1176_5.INIT1 = 16'hf555;
    defparam add_1176_5.INJECT1_0 = "NO";
    defparam add_1176_5.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_19 (.A0(multOut[17]), .B0(n16618), .C0(addOut[17]), 
          .D0(addIn2_28__N_1207[17]), .A1(multOut[18]), .B1(n16618), .C1(addOut[18]), 
          .D1(addIn2_28__N_1207[18]), .CIN(n18565), .COUT(n18566), .S0(n121[17]), 
          .S1(n121[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_19.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_19.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_19.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_19.INJECT1_1 = "NO";
    LUT4 mux_1800_i4_3_lut_4_lut (.A(ss[2]), .B(n21553), .C(\speed_m1[3] ), 
         .D(subIn2_24__N_1301[3]), .Z(subIn2_24__N_1114[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_1800_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut_adj_71 (.A(n22208), .B(n920), .C(addOut[15]), 
         .D(n3635), .Z(intgOut0_28__N_735[15])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_71.init = 16'h1110;
    CCU2D add_191_5 (.A0(Out3[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18440), 
          .COUT(n18441), .S0(n1208[3]), .S1(n1208[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_5.INIT0 = 16'h5aaa;
    defparam add_191_5.INIT1 = 16'h5aaa;
    defparam add_191_5.INJECT1_0 = "NO";
    defparam add_191_5.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_17 (.A0(multOut[15]), .B0(n16618), .C0(addOut[15]), 
          .D0(addIn2_28__N_1207[15]), .A1(multOut[16]), .B1(n16618), .C1(addOut[16]), 
          .D1(addIn2_28__N_1207[16]), .CIN(n18564), .COUT(n18565), .S0(n121[15]), 
          .S1(n121[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_17.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_17.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_17.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_17.INJECT1_1 = "NO";
    CCU2D add_15799_15 (.A0(addOut[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18699), .COUT(n18700));
    defparam add_15799_15.INIT0 = 16'hf555;
    defparam add_15799_15.INIT1 = 16'h0aaa;
    defparam add_15799_15.INJECT1_0 = "NO";
    defparam add_15799_15.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_15 (.A0(multOut[13]), .B0(n16618), .C0(addOut[13]), 
          .D0(addIn2_28__N_1207[13]), .A1(multOut[14]), .B1(n16618), .C1(addOut[14]), 
          .D1(addIn2_28__N_1207[14]), .CIN(n18563), .COUT(n18564), .S0(n121[13]), 
          .S1(n121[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_15.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_15.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_15.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_15.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i24 (.BLUT(n618[23]), .ALUT(addIn2_28__N_1337[23]), 
          .C0(n20447), .Z(addIn2_28__N_1207[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D addOut_2063_add_4_13 (.A0(multOut[11]), .B0(n16618), .C0(addOut[11]), 
          .D0(addIn2_28__N_1207[11]), .A1(multOut[12]), .B1(n16618), .C1(addOut[12]), 
          .D1(addIn2_28__N_1207[12]), .CIN(n18562), .COUT(n18563), .S0(n121[11]), 
          .S1(n121[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_13.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_13.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_13.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_13.INJECT1_1 = "NO";
    CCU2D add_15799_13 (.A0(addOut[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18698), .COUT(n18699));
    defparam add_15799_13.INIT0 = 16'h0aaa;
    defparam add_15799_13.INIT1 = 16'h0aaa;
    defparam add_15799_13.INJECT1_0 = "NO";
    defparam add_15799_13.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i23 (.BLUT(n618[22]), .ALUT(addIn2_28__N_1337[22]), 
          .C0(n20447), .Z(addIn2_28__N_1207[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1176_3 (.A0(n1208[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18512), 
          .COUT(n18513), .S0(n2188[1]), .S1(n2188[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(351[20:29])
    defparam add_1176_3.INIT0 = 16'hf555;
    defparam add_1176_3.INIT1 = 16'hf555;
    defparam add_1176_3.INJECT1_0 = "NO";
    defparam add_1176_3.INJECT1_1 = "NO";
    CCU2D add_15799_11 (.A0(addOut[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18697), .COUT(n18698));
    defparam add_15799_11.INIT0 = 16'h0aaa;
    defparam add_15799_11.INIT1 = 16'h0aaa;
    defparam add_15799_11.INJECT1_0 = "NO";
    defparam add_15799_11.INJECT1_1 = "NO";
    CCU2D add_191_3 (.A0(Out3[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18439), 
          .COUT(n18440), .S0(n1208[1]), .S1(n1208[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_3.INIT0 = 16'h5aaa;
    defparam add_191_3.INIT1 = 16'h5aaa;
    defparam add_191_3.INJECT1_0 = "NO";
    defparam add_191_3.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_11 (.A0(multOut[9]), .B0(n16618), .C0(addOut[9]), 
          .D0(addIn2_28__N_1207[9]), .A1(multOut[10]), .B1(n16618), .C1(addOut[10]), 
          .D1(addIn2_28__N_1207[10]), .CIN(n18561), .COUT(n18562), .S0(n121[9]), 
          .S1(n121[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_11.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_11.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_11.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_11.INJECT1_1 = "NO";
    CCU2D add_191_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[13]), .B1(n18859), .C1(n18860), .D1(Out3[28]), .COUT(n18439), 
          .S1(n1208[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_1.INIT0 = 16'hF000;
    defparam add_191_1.INIT1 = 16'h56aa;
    defparam add_191_1.INJECT1_0 = "NO";
    defparam add_191_1.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i22 (.BLUT(n618[21]), .ALUT(addIn2_28__N_1337[21]), 
          .C0(n20447), .Z(addIn2_28__N_1207[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1176_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1208[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18512), 
          .S1(n2188[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(351[20:29])
    defparam add_1176_1.INIT0 = 16'hF000;
    defparam add_1176_1.INIT1 = 16'h0aaa;
    defparam add_1176_1.INJECT1_0 = "NO";
    defparam add_1176_1.INJECT1_1 = "NO";
    CCU2D add_15799_9 (.A0(addOut[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18696), .COUT(n18697));
    defparam add_15799_9.INIT0 = 16'h0aaa;
    defparam add_15799_9.INIT1 = 16'hf555;
    defparam add_15799_9.INJECT1_0 = "NO";
    defparam add_15799_9.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_9 (.A0(multOut[7]), .B0(n16618), .C0(addOut[7]), 
          .D0(addIn2_28__N_1207[7]), .A1(multOut[8]), .B1(n16618), .C1(addOut[8]), 
          .D1(addIn2_28__N_1207[8]), .CIN(n18560), .COUT(n18561), .S0(n121[7]), 
          .S1(n121[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_9.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_9.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_9.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_282_3_lut_4_lut_4_lut (.A(n21554), .B(n21530), .C(n35), 
         .D(n21552), .Z(n21491)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i1_2_lut_rep_282_3_lut_4_lut_4_lut.init = 16'hc0d0;
    CCU2D add_15799_7 (.A0(addOut[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18695), .COUT(n18696));
    defparam add_15799_7.INIT0 = 16'h0aaa;
    defparam add_15799_7.INIT1 = 16'h0aaa;
    defparam add_15799_7.INJECT1_0 = "NO";
    defparam add_15799_7.INJECT1_1 = "NO";
    CCU2D add_15799_5 (.A0(addOut[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18694), .COUT(n18695));
    defparam add_15799_5.INIT0 = 16'hf555;
    defparam add_15799_5.INIT1 = 16'hf555;
    defparam add_15799_5.INJECT1_0 = "NO";
    defparam add_15799_5.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_7 (.A0(multOut[5]), .B0(n16618), .C0(addOut[5]), 
          .D0(addIn2_28__N_1207[5]), .A1(multOut[6]), .B1(n16618), .C1(addOut[6]), 
          .D1(addIn2_28__N_1207[6]), .CIN(n18559), .COUT(n18560), .S0(n121[5]), 
          .S1(n121[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_7.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_7.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_7.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_7.INJECT1_1 = "NO";
    CCU2D add_1175_11 (.A0(n1187[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18511), 
          .S0(n2176[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(343[20:29])
    defparam add_1175_11.INIT0 = 16'hf555;
    defparam add_1175_11.INIT1 = 16'h0000;
    defparam add_1175_11.INJECT1_0 = "NO";
    defparam add_1175_11.INJECT1_1 = "NO";
    CCU2D add_1175_9 (.A0(n1187[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18510), 
          .COUT(n18511), .S0(n2176[7]), .S1(n2176[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(343[20:29])
    defparam add_1175_9.INIT0 = 16'hf555;
    defparam add_1175_9.INIT1 = 16'hf555;
    defparam add_1175_9.INJECT1_0 = "NO";
    defparam add_1175_9.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_5 (.A0(multOut[3]), .B0(n16618), .C0(addOut[3]), 
          .D0(addIn2_28__N_1207[3]), .A1(multOut[4]), .B1(n16618), .C1(addOut[4]), 
          .D1(addIn2_28__N_1207[4]), .CIN(n18558), .COUT(n18559), .S0(n121[3]), 
          .S1(n121[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_5.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_5.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_5.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_5.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_3 (.A0(multOut[1]), .B0(n16618), .C0(addOut[1]), 
          .D0(addIn2_28__N_1207[1]), .A1(multOut[2]), .B1(n16618), .C1(addOut[2]), 
          .D1(addIn2_28__N_1207[2]), .CIN(n18557), .COUT(n18558), .S0(n121[1]), 
          .S1(n121[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_3.INIT0 = 16'h569a;
    defparam addOut_2063_add_4_3.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_3.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_3.INJECT1_1 = "NO";
    CCU2D add_1175_7 (.A0(n1187[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18509), 
          .COUT(n18510), .S0(n2176[5]), .S1(n2176[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(343[20:29])
    defparam add_1175_7.INIT0 = 16'hf555;
    defparam add_1175_7.INIT1 = 16'hf555;
    defparam add_1175_7.INJECT1_0 = "NO";
    defparam add_1175_7.INJECT1_1 = "NO";
    CCU2D addOut_2063_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(multOut[0]), .B1(n16618), .C1(addOut[0]), 
          .D1(addIn2_28__N_1207[0]), .COUT(n18557), .S1(n121[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063_add_4_1.INIT0 = 16'hF000;
    defparam addOut_2063_add_4_1.INIT1 = 16'h569a;
    defparam addOut_2063_add_4_1.INJECT1_0 = "NO";
    defparam addOut_2063_add_4_1.INJECT1_1 = "NO";
    CCU2D add_187_17 (.A0(Out2[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18438), 
          .S0(n1187[15]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_17.INIT0 = 16'h5aaa;
    defparam add_187_17.INIT1 = 16'h0000;
    defparam add_187_17.INJECT1_0 = "NO";
    defparam add_187_17.INJECT1_1 = "NO";
    CCU2D add_187_15 (.A0(Out2[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18437), 
          .COUT(n18438), .S0(n1187[13]), .S1(n1187[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_15.INIT0 = 16'h5aaa;
    defparam add_187_15.INIT1 = 16'h5aaa;
    defparam add_187_15.INJECT1_0 = "NO";
    defparam add_187_15.INJECT1_1 = "NO";
    CCU2D add_15799_3 (.A0(addOut[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18693), .COUT(n18694));
    defparam add_15799_3.INIT0 = 16'hf555;
    defparam add_15799_3.INIT1 = 16'hf555;
    defparam add_15799_3.INJECT1_0 = "NO";
    defparam add_15799_3.INJECT1_1 = "NO";
    CCU2D add_15799_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[0]), .B1(addOut[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18693));
    defparam add_15799_1.INIT0 = 16'hF000;
    defparam add_15799_1.INIT1 = 16'ha666;
    defparam add_15799_1.INJECT1_0 = "NO";
    defparam add_15799_1.INJECT1_1 = "NO";
    CCU2D add_15800_21 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18692), .S1(n56));
    defparam add_15800_21.INIT0 = 16'h5555;
    defparam add_15800_21.INIT1 = 16'h0000;
    defparam add_15800_21.INJECT1_0 = "NO";
    defparam add_15800_21.INJECT1_1 = "NO";
    CCU2D add_15800_19 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18691), .COUT(n18692));
    defparam add_15800_19.INIT0 = 16'hf555;
    defparam add_15800_19.INIT1 = 16'hf555;
    defparam add_15800_19.INJECT1_0 = "NO";
    defparam add_15800_19.INJECT1_1 = "NO";
    CCU2D add_15800_17 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18690), .COUT(n18691));
    defparam add_15800_17.INIT0 = 16'hf555;
    defparam add_15800_17.INIT1 = 16'hf555;
    defparam add_15800_17.INJECT1_0 = "NO";
    defparam add_15800_17.INJECT1_1 = "NO";
    CCU2D add_1175_5 (.A0(n1187[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18508), 
          .COUT(n18509), .S0(n2176[3]), .S1(n2176[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(343[20:29])
    defparam add_1175_5.INIT0 = 16'hf555;
    defparam add_1175_5.INIT1 = 16'hf555;
    defparam add_1175_5.INJECT1_0 = "NO";
    defparam add_1175_5.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i21 (.BLUT(n618[20]), .ALUT(addIn2_28__N_1337[20]), 
          .C0(n20447), .Z(addIn2_28__N_1207[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i14128_2_lut_rep_390 (.A(ss[1]), .B(ss[3]), .Z(n21599)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14128_2_lut_rep_390.init = 16'heeee;
    CCU2D add_1175_3 (.A0(n1187[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18507), 
          .COUT(n18508), .S0(n2176[1]), .S1(n2176[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(343[20:29])
    defparam add_1175_3.INIT0 = 16'hf555;
    defparam add_1175_3.INIT1 = 16'hf555;
    defparam add_1175_3.INJECT1_0 = "NO";
    defparam add_1175_3.INJECT1_1 = "NO";
    LUT4 i17838_2_lut_rep_278_2_lut_3_lut_4_lut_4_lut (.A(n21554), .B(n21530), 
         .C(n35), .D(n21552), .Z(n21487)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B (C+(D))))) */ ;
    defparam i17838_2_lut_rep_278_2_lut_3_lut_4_lut_4_lut.init = 16'h0c0d;
    CCU2D add_187_13 (.A0(Out2[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18436), 
          .COUT(n18437), .S0(n1187[11]), .S1(n1187[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_13.INIT0 = 16'h5aaa;
    defparam add_187_13.INIT1 = 16'h5aaa;
    defparam add_187_13.INJECT1_0 = "NO";
    defparam add_187_13.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut (.A(ss[1]), .B(ss[3]), .C(n22199), .D(ss[0]), 
         .Z(n18815)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_187_11 (.A0(Out2[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18435), 
          .COUT(n18436), .S0(n1187[9]), .S1(n1187[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_11.INIT0 = 16'h5aaa;
    defparam add_187_11.INIT1 = 16'h5aaa;
    defparam add_187_11.INJECT1_0 = "NO";
    defparam add_187_11.INJECT1_1 = "NO";
    CCU2D add_15800_15 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18689), .COUT(n18690));
    defparam add_15800_15.INIT0 = 16'hf555;
    defparam add_15800_15.INIT1 = 16'hf555;
    defparam add_15800_15.INJECT1_0 = "NO";
    defparam add_15800_15.INJECT1_1 = "NO";
    CCU2D add_1175_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1187[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18507), 
          .S1(n2176[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(343[20:29])
    defparam add_1175_1.INIT0 = 16'hF000;
    defparam add_1175_1.INIT1 = 16'h0aaa;
    defparam add_1175_1.INJECT1_0 = "NO";
    defparam add_1175_1.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i20 (.BLUT(n618[19]), .ALUT(addIn2_28__N_1337[19]), 
          .C0(n20447), .Z(addIn2_28__N_1207[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_137_i1_3_lut_4_lut_4_lut (.A(n21554), .B(n588[0]), .C(intgOut3[0]), 
         .D(n21552), .Z(n618[0])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i1_3_lut_4_lut_4_lut.init = 16'hccd8;
    FD1P3IX dutyout_m2_i0_i0 (.D(n2164[0]), .SP(clk_N_683_enable_392), .CD(n12648), 
            .CK(clk_N_683), .Q(PWMdut_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i0.GSR = "DISABLED";
    LUT4 mux_137_i17_3_lut_4_lut_4_lut (.A(n21554), .B(n588[16]), .C(intgOut3[16]), 
         .D(n21552), .Z(n618[16])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i17_3_lut_4_lut_4_lut.init = 16'hccd8;
    FD1P3IX dutyout_m1_i0_i0 (.D(n2152[0]), .SP(clk_N_683_enable_392), .CD(n12639), 
            .CK(clk_N_683), .Q(PWMdut_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i0.GSR = "DISABLED";
    LUT4 mux_137_i16_3_lut_4_lut_4_lut (.A(n21554), .B(n588[15]), .C(intgOut3[15]), 
         .D(n21552), .Z(n618[15])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i16_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i15_3_lut_4_lut_4_lut (.A(n21554), .B(n588[14]), .C(intgOut3[14]), 
         .D(n21552), .Z(n618[14])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i15_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i14_3_lut_4_lut_4_lut (.A(n21554), .B(n588[13]), .C(intgOut3[13]), 
         .D(n21552), .Z(n618[13])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX addIn2_28__I_29_i19 (.BLUT(n618[18]), .ALUT(addIn2_28__N_1337[18]), 
          .C0(n20447), .Z(addIn2_28__N_1207[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1_2_lut_3_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n19668)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_392 (.A(ss[0]), .B(ss[3]), .Z(n21601)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_392.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_72 (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n19776)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_3_lut_adj_72.init = 16'hfbfb;
    LUT4 mux_137_i13_3_lut_4_lut_4_lut (.A(n21554), .B(n588[12]), .C(intgOut3[12]), 
         .D(n21552), .Z(n618[12])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i13_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i12_3_lut_4_lut_4_lut (.A(n21554), .B(n588[11]), .C(intgOut3[11]), 
         .D(n21552), .Z(n618[11])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i11_3_lut_4_lut_4_lut (.A(n21554), .B(n588[10]), .C(intgOut3[10]), 
         .D(n21552), .Z(n618[10])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i10_3_lut_4_lut_4_lut (.A(n21554), .B(n588[9]), .C(intgOut3[9]), 
         .D(n21552), .Z(n618[9])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i10_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX addIn2_28__I_29_i18 (.BLUT(n618[17]), .ALUT(addIn2_28__N_1337[17]), 
          .C0(n20447), .Z(addIn2_28__N_1207[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    FD1P3IX dutyout_m2_i0_i1 (.D(n2164[1]), .SP(clk_N_683_enable_392), .CD(n12648), 
            .CK(clk_N_683), .Q(PWMdut_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i1.GSR = "DISABLED";
    LUT4 mux_137_i2_3_lut_4_lut_4_lut (.A(n21554), .B(n588[1]), .C(intgOut3[1]), 
         .D(n21552), .Z(n618[1])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i2_3_lut_4_lut_4_lut.init = 16'hccd8;
    CCU2D add_15800_13 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18688), .COUT(n18689));
    defparam add_15800_13.INIT0 = 16'hf555;
    defparam add_15800_13.INIT1 = 16'hf555;
    defparam add_15800_13.INJECT1_0 = "NO";
    defparam add_15800_13.INJECT1_1 = "NO";
    CCU2D add_1174_11 (.A0(n1166[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18506), 
          .S0(n2164[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(335[20:29])
    defparam add_1174_11.INIT0 = 16'hf555;
    defparam add_1174_11.INIT1 = 16'h0000;
    defparam add_1174_11.INJECT1_0 = "NO";
    defparam add_1174_11.INJECT1_1 = "NO";
    CCU2D add_187_9 (.A0(Out2[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18434), 
          .COUT(n18435), .S0(n1187[7]), .S1(n1187[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_9.INIT0 = 16'h5aaa;
    defparam add_187_9.INIT1 = 16'h5aaa;
    defparam add_187_9.INJECT1_0 = "NO";
    defparam add_187_9.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i9 (.BLUT(n618[8]), .ALUT(addIn2_28__N_1337[8]), 
          .C0(n20447), .Z(addIn2_28__N_1207[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_15800_11 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18687), .COUT(n18688));
    defparam add_15800_11.INIT0 = 16'hf555;
    defparam add_15800_11.INIT1 = 16'hf555;
    defparam add_15800_11.INJECT1_0 = "NO";
    defparam add_15800_11.INJECT1_1 = "NO";
    CCU2D add_15800_9 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18686), .COUT(n18687));
    defparam add_15800_9.INIT0 = 16'hf555;
    defparam add_15800_9.INIT1 = 16'hf555;
    defparam add_15800_9.INJECT1_0 = "NO";
    defparam add_15800_9.INJECT1_1 = "NO";
    CCU2D add_15800_7 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18685), .COUT(n18686));
    defparam add_15800_7.INIT0 = 16'hf555;
    defparam add_15800_7.INIT1 = 16'hf555;
    defparam add_15800_7.INJECT1_0 = "NO";
    defparam add_15800_7.INJECT1_1 = "NO";
    CCU2D add_187_7 (.A0(Out2[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18433), 
          .COUT(n18434), .S0(n1187[5]), .S1(n1187[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_7.INIT0 = 16'h5aaa;
    defparam add_187_7.INIT1 = 16'h5aaa;
    defparam add_187_7.INJECT1_0 = "NO";
    defparam add_187_7.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i7 (.BLUT(n618[6]), .ALUT(addIn2_28__N_1337[6]), 
          .C0(n20447), .Z(addIn2_28__N_1207[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1174_9 (.A0(n1166[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18505), 
          .COUT(n18506), .S0(n2164[7]), .S1(n2164[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(335[20:29])
    defparam add_1174_9.INIT0 = 16'hf555;
    defparam add_1174_9.INIT1 = 16'hf555;
    defparam add_1174_9.INJECT1_0 = "NO";
    defparam add_1174_9.INJECT1_1 = "NO";
    CCU2D add_15800_5 (.A0(speed_set_m4[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18684), .COUT(n18685));
    defparam add_15800_5.INIT0 = 16'hf555;
    defparam add_15800_5.INIT1 = 16'hf555;
    defparam add_15800_5.INJECT1_0 = "NO";
    defparam add_15800_5.INJECT1_1 = "NO";
    CCU2D add_1174_7 (.A0(n1166[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18504), 
          .COUT(n18505), .S0(n2164[5]), .S1(n2164[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(335[20:29])
    defparam add_1174_7.INIT0 = 16'hf555;
    defparam add_1174_7.INIT1 = 16'hf555;
    defparam add_1174_7.INJECT1_0 = "NO";
    defparam add_1174_7.INJECT1_1 = "NO";
    CCU2D add_15800_3 (.A0(speed_set_m4[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18683), .COUT(n18684));
    defparam add_15800_3.INIT0 = 16'hf555;
    defparam add_15800_3.INIT1 = 16'hf555;
    defparam add_15800_3.INJECT1_0 = "NO";
    defparam add_15800_3.INJECT1_1 = "NO";
    CCU2D add_187_5 (.A0(Out2[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18432), 
          .COUT(n18433), .S0(n1187[3]), .S1(n1187[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_5.INIT0 = 16'h5aaa;
    defparam add_187_5.INIT1 = 16'h5aaa;
    defparam add_187_5.INJECT1_0 = "NO";
    defparam add_187_5.INJECT1_1 = "NO";
    CCU2D add_187_3 (.A0(Out2[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18431), 
          .COUT(n18432), .S0(n1187[1]), .S1(n1187[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_3.INIT0 = 16'h5aaa;
    defparam add_187_3.INIT1 = 16'h5aaa;
    defparam add_187_3.INJECT1_0 = "NO";
    defparam add_187_3.INJECT1_1 = "NO";
    CCU2D add_15800_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[0]), .B1(speed_set_m4[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18683));
    defparam add_15800_1.INIT0 = 16'hF000;
    defparam add_15800_1.INIT1 = 16'ha666;
    defparam add_15800_1.INJECT1_0 = "NO";
    defparam add_15800_1.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i3 (.BLUT(n618[2]), .ALUT(addIn2_28__N_1337[2]), 
          .C0(n20447), .Z(addIn2_28__N_1207[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_1174_5 (.A0(n1166[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18503), 
          .COUT(n18504), .S0(n2164[3]), .S1(n2164[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(335[20:29])
    defparam add_1174_5.INIT0 = 16'hf555;
    defparam add_1174_5.INIT1 = 16'hf555;
    defparam add_1174_5.INJECT1_0 = "NO";
    defparam add_1174_5.INJECT1_1 = "NO";
    CCU2D add_1174_3 (.A0(n1166[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18502), 
          .COUT(n18503), .S0(n2164[1]), .S1(n2164[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(335[20:29])
    defparam add_1174_3.INIT0 = 16'hf555;
    defparam add_1174_3.INIT1 = 16'hf555;
    defparam add_1174_3.INJECT1_0 = "NO";
    defparam add_1174_3.INJECT1_1 = "NO";
    CCU2D add_1174_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1166[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18502), 
          .S1(n2164[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(335[20:29])
    defparam add_1174_1.INIT0 = 16'hF000;
    defparam add_1174_1.INIT1 = 16'h0aaa;
    defparam add_1174_1.INJECT1_0 = "NO";
    defparam add_1174_1.INJECT1_1 = "NO";
    CCU2D add_187_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[13]), .B1(n18862), .C1(n18863), .D1(Out2[28]), .COUT(n18431), 
          .S1(n1187[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(316[17:21])
    defparam add_187_1.INIT0 = 16'hF000;
    defparam add_187_1.INIT1 = 16'h56aa;
    defparam add_187_1.INJECT1_0 = "NO";
    defparam add_187_1.INJECT1_1 = "NO";
    CCU2D add_183_17 (.A0(Out1[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18430), 
          .S0(n1166[15]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_17.INIT0 = 16'h5aaa;
    defparam add_183_17.INIT1 = 16'h0000;
    defparam add_183_17.INJECT1_0 = "NO";
    defparam add_183_17.INJECT1_1 = "NO";
    CCU2D sub_16_rep_2_add_2_25 (.A0(n16636), .B0(n16636), .C0(n27[21]), 
          .D0(n2244[21]), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18501), .S0(subOut_24__N_1135[24]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_25.INIT0 = 16'h569a;
    defparam sub_16_rep_2_add_2_25.INIT1 = 16'h0000;
    defparam sub_16_rep_2_add_2_25.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_25.INJECT1_1 = "NO";
    CCU2D add_183_15 (.A0(Out1[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18429), 
          .COUT(n18430), .S0(n1166[13]), .S1(n1166[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_15.INIT0 = 16'h5aaa;
    defparam add_183_15.INIT1 = 16'h5aaa;
    defparam add_183_15.INJECT1_0 = "NO";
    defparam add_183_15.INJECT1_1 = "NO";
    CCU2D add_15801_21 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18682), .S1(n49));
    defparam add_15801_21.INIT0 = 16'h5555;
    defparam add_15801_21.INIT1 = 16'h0000;
    defparam add_15801_21.INJECT1_0 = "NO";
    defparam add_15801_21.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i8 (.BLUT(n618[7]), .ALUT(addIn2_28__N_1337[7]), 
          .C0(n20447), .Z(addIn2_28__N_1207[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_15801_19 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18681), .COUT(n18682));
    defparam add_15801_19.INIT0 = 16'hf555;
    defparam add_15801_19.INIT1 = 16'hf555;
    defparam add_15801_19.INJECT1_0 = "NO";
    defparam add_15801_19.INJECT1_1 = "NO";
    CCU2D add_15801_17 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18680), .COUT(n18681));
    defparam add_15801_17.INIT0 = 16'hf555;
    defparam add_15801_17.INIT1 = 16'hf555;
    defparam add_15801_17.INJECT1_0 = "NO";
    defparam add_15801_17.INJECT1_1 = "NO";
    CCU2D add_15801_15 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18679), .COUT(n18680));
    defparam add_15801_15.INIT0 = 16'hf555;
    defparam add_15801_15.INIT1 = 16'hf555;
    defparam add_15801_15.INJECT1_0 = "NO";
    defparam add_15801_15.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i4 (.BLUT(n618[3]), .ALUT(addIn2_28__N_1337[3]), 
          .C0(n20447), .Z(addIn2_28__N_1207[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_183_13 (.A0(Out1[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18428), 
          .COUT(n18429), .S0(n1166[11]), .S1(n1166[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_13.INIT0 = 16'h5aaa;
    defparam add_183_13.INIT1 = 16'h5aaa;
    defparam add_183_13.INJECT1_0 = "NO";
    defparam add_183_13.INJECT1_1 = "NO";
    CCU2D add_183_11 (.A0(Out1[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18427), 
          .COUT(n18428), .S0(n1166[9]), .S1(n1166[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_11.INIT0 = 16'h5aaa;
    defparam add_183_11.INIT1 = 16'h5aaa;
    defparam add_183_11.INJECT1_0 = "NO";
    defparam add_183_11.INJECT1_1 = "NO";
    CCU2D add_15801_13 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18678), .COUT(n18679));
    defparam add_15801_13.INIT0 = 16'hf555;
    defparam add_15801_13.INIT1 = 16'hf555;
    defparam add_15801_13.INJECT1_0 = "NO";
    defparam add_15801_13.INJECT1_1 = "NO";
    CCU2D add_15801_11 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18677), .COUT(n18678));
    defparam add_15801_11.INIT0 = 16'hf555;
    defparam add_15801_11.INIT1 = 16'hf555;
    defparam add_15801_11.INJECT1_0 = "NO";
    defparam add_15801_11.INJECT1_1 = "NO";
    CCU2D sub_16_rep_2_add_2_23 (.A0(n16636), .B0(n16636), .C0(n27[20]), 
          .D0(n2244[20]), .A1(n16636), .B1(n16636), .C1(n27[21]), .D1(n2244[21]), 
          .CIN(n18500), .COUT(n18501), .S0(subOut_24__N_1135[20]), .S1(subOut_24__N_1135[21]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_23.INIT0 = 16'h569a;
    defparam sub_16_rep_2_add_2_23.INIT1 = 16'h569a;
    defparam sub_16_rep_2_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_16_rep_2_add_2_21 (.A0(subIn2[18]), .B0(n16636), .C0(n27[18]), 
          .D0(n2244[18]), .A1(n7), .B1(n16636), .C1(n27[19]), .D1(n2244[19]), 
          .CIN(n18499), .COUT(n18500), .S0(subOut_24__N_1135[18]), .S1(subOut_24__N_1135[19]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_21.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_21.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_16_rep_2_add_2_19 (.A0(subIn2[16]), .B0(n16636), .C0(n27[16]), 
          .D0(n2244[16]), .A1(subIn2[17]), .B1(n16636), .C1(n27[17]), 
          .D1(n2244[17]), .CIN(n18498), .COUT(n18499), .S0(subOut_24__N_1135[16]), 
          .S1(subOut_24__N_1135[17]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_19.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_19.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_19.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i5 (.BLUT(n618[4]), .ALUT(addIn2_28__N_1337[4]), 
          .C0(n20447), .Z(addIn2_28__N_1207[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1_2_lut_rep_398 (.A(n22199), .B(ss[1]), .Z(n21607)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_398.init = 16'heeee;
    CCU2D add_183_9 (.A0(Out1[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18426), 
          .COUT(n18427), .S0(n1166[7]), .S1(n1166[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_9.INIT0 = 16'h5aaa;
    defparam add_183_9.INIT1 = 16'h5aaa;
    defparam add_183_9.INJECT1_0 = "NO";
    defparam add_183_9.INJECT1_1 = "NO";
    CCU2D add_183_7 (.A0(Out1[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18425), 
          .COUT(n18426), .S0(n1166[5]), .S1(n1166[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_7.INIT0 = 16'h5aaa;
    defparam add_183_7.INIT1 = 16'h5aaa;
    defparam add_183_7.INJECT1_0 = "NO";
    defparam add_183_7.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i6 (.BLUT(n618[5]), .ALUT(addIn2_28__N_1337[5]), 
          .C0(n20447), .Z(addIn2_28__N_1207[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D sub_16_rep_2_add_2_17 (.A0(subIn2[14]), .B0(n16636), .C0(n27[14]), 
          .D0(n2244[14]), .A1(subIn2[15]), .B1(n16636), .C1(n27[15]), 
          .D1(n2244[15]), .CIN(n18497), .COUT(n18498), .S0(subOut_24__N_1135[14]), 
          .S1(subOut_24__N_1135[15]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_17.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_17.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_17.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i2 (.BLUT(n618[1]), .ALUT(addIn2_28__N_1337[1]), 
          .C0(n20447), .Z(addIn2_28__N_1207[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D sub_16_rep_2_add_2_15 (.A0(subIn2[12]), .B0(n16636), .C0(n27[12]), 
          .D0(n2244[12]), .A1(subIn2[13]), .B1(n16636), .C1(n27[13]), 
          .D1(n2244[13]), .CIN(n18496), .COUT(n18497), .S0(subOut_24__N_1135[12]), 
          .S1(subOut_24__N_1135[13]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_15.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_15.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_15.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_339_4_lut (.A(ss[2]), .B(ss[1]), .C(ss[3]), .D(n22208), 
         .Z(n21548)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i1_3_lut_rep_339_4_lut.init = 16'h001e;
    LUT4 mux_137_i6_3_lut_4_lut_4_lut (.A(n21554), .B(n588[5]), .C(intgOut3[5]), 
         .D(n21552), .Z(n618[5])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i6_3_lut_4_lut_4_lut.init = 16'hccd8;
    CCU2D sub_16_rep_2_add_2_13 (.A0(subIn2[10]), .B0(n16636), .C0(n27[10]), 
          .D0(n2244[10]), .A1(subIn2[11]), .B1(n16636), .C1(n27[11]), 
          .D1(n2244[11]), .CIN(n18495), .COUT(n18496), .S0(subOut_24__N_1135[10]), 
          .S1(subOut_24__N_1135[11]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_13.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_13.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_399 (.A(ss[0]), .B(ss[3]), .Z(n21608)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_399.init = 16'heeee;
    CCU2D add_183_5 (.A0(Out1[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18424), 
          .COUT(n18425), .S0(n1166[3]), .S1(n1166[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_5.INIT0 = 16'h5aaa;
    defparam add_183_5.INIT1 = 16'h5aaa;
    defparam add_183_5.INJECT1_0 = "NO";
    defparam add_183_5.INJECT1_1 = "NO";
    LUT4 i2_2_lut_rep_360_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), 
         .D(ss[2]), .Z(n21569)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i2_2_lut_rep_360_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_183_3 (.A0(Out1[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18423), 
          .COUT(n18424), .S0(n1166[1]), .S1(n1166[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_3.INIT0 = 16'h5aaa;
    defparam add_183_3.INIT1 = 16'h5aaa;
    defparam add_183_3.INJECT1_0 = "NO";
    defparam add_183_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_73 (.A(n22208), .B(n920), .C(addOut[20]), 
         .D(n3635), .Z(intgOut0_28__N_735[20])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_73.init = 16'h1110;
    LUT4 mux_137_i5_3_lut_4_lut_4_lut (.A(n21554), .B(n588[4]), .C(intgOut3[4]), 
         .D(n21552), .Z(n618[4])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i5_3_lut_4_lut_4_lut.init = 16'hccd8;
    CCU2D add_15801_9 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18676), .COUT(n18677));
    defparam add_15801_9.INIT0 = 16'hf555;
    defparam add_15801_9.INIT1 = 16'hf555;
    defparam add_15801_9.INJECT1_0 = "NO";
    defparam add_15801_9.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i10 (.BLUT(n618[9]), .ALUT(addIn2_28__N_1337[9]), 
          .C0(n20447), .Z(addIn2_28__N_1207[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 i1_3_lut_4_lut_adj_74 (.A(n22208), .B(n920), .C(addOut[21]), 
         .D(n3635), .Z(intgOut0_28__N_735[21])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_74.init = 16'h1110;
    LUT4 mux_137_i4_3_lut_4_lut_4_lut (.A(n21554), .B(n588[3]), .C(intgOut3[3]), 
         .D(n21552), .Z(n618[3])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i4_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i1_3_lut_4_lut_adj_75 (.A(n22208), .B(n920), .C(addOut[22]), 
         .D(n3635), .Z(intgOut0_28__N_735[22])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_75.init = 16'h1110;
    CCU2D add_183_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[13]), .B1(n18821), .C1(n18822), .D1(Out1[28]), .COUT(n18423), 
          .S1(n1166[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(315[17:21])
    defparam add_183_1.INIT0 = 16'hF000;
    defparam add_183_1.INIT1 = 16'h56aa;
    defparam add_183_1.INJECT1_0 = "NO";
    defparam add_183_1.INJECT1_1 = "NO";
    CCU2D add_15801_7 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18675), .COUT(n18676));
    defparam add_15801_7.INIT0 = 16'hf555;
    defparam add_15801_7.INIT1 = 16'hf555;
    defparam add_15801_7.INJECT1_0 = "NO";
    defparam add_15801_7.INJECT1_1 = "NO";
    CCU2D add_15801_5 (.A0(speed_set_m3[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18674), .COUT(n18675));
    defparam add_15801_5.INIT0 = 16'hf555;
    defparam add_15801_5.INIT1 = 16'hf555;
    defparam add_15801_5.INJECT1_0 = "NO";
    defparam add_15801_5.INJECT1_1 = "NO";
    CCU2D sub_16_rep_2_add_2_11 (.A0(subIn2[8]), .B0(n16636), .C0(n27[8]), 
          .D0(n2244[8]), .A1(subIn2[9]), .B1(n16636), .C1(n27[9]), .D1(n2244[9]), 
          .CIN(n18494), .COUT(n18495), .S0(subOut_24__N_1135[8]), .S1(subOut_24__N_1135[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_11.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_11.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_11.INJECT1_1 = "NO";
    PFUMX addIn2_28__I_29_i11 (.BLUT(n618[10]), .ALUT(addIn2_28__N_1337[10]), 
          .C0(n20447), .Z(addIn2_28__N_1207[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_137_i8_3_lut_4_lut_4_lut (.A(n21554), .B(n588[7]), .C(intgOut3[7]), 
         .D(n21552), .Z(n618[7])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i8_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i3_3_lut_4_lut_4_lut (.A(n21554), .B(n588[2]), .C(intgOut3[2]), 
         .D(n21552), .Z(n618[2])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i3_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i7_3_lut_4_lut_4_lut (.A(n21554), .B(n588[6]), .C(intgOut3[6]), 
         .D(n21552), .Z(n618[6])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i7_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i9_3_lut_4_lut_4_lut (.A(n21554), .B(n588[8]), .C(intgOut3[8]), 
         .D(n21552), .Z(n618[8])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i9_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX i18138 (.BLUT(n21609), .ALUT(n21610), .C0(n22208), .Z(clk_N_683_enable_241));
    LUT4 mux_137_i18_3_lut_4_lut_4_lut (.A(n21554), .B(n588[17]), .C(intgOut3[17]), 
         .D(n21552), .Z(n618[17])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i18_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i19_3_lut_4_lut_4_lut (.A(n21554), .B(n588[18]), .C(intgOut3[18]), 
         .D(n21552), .Z(n618[18])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i19_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i20_3_lut_4_lut_4_lut (.A(n21554), .B(n588[19]), .C(intgOut3[19]), 
         .D(n21552), .Z(n618[19])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i20_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX addIn2_28__I_29_i12 (.BLUT(n618[11]), .ALUT(addIn2_28__N_1337[11]), 
          .C0(n20447), .Z(addIn2_28__N_1207[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_137_i21_3_lut_4_lut_4_lut (.A(n21554), .B(n588[20]), .C(intgOut3[20]), 
         .D(n21552), .Z(n618[20])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i21_3_lut_4_lut_4_lut.init = 16'hccd8;
    CCU2D add_179_17 (.A0(Out0[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18422), 
          .S0(n1145[15]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_17.INIT0 = 16'h5aaa;
    defparam add_179_17.INIT1 = 16'h0000;
    defparam add_179_17.INJECT1_0 = "NO";
    defparam add_179_17.INJECT1_1 = "NO";
    FD1S3AY ss_i4_rep_411 (.D(n19725), .CK(clk_N_683), .Q(n22208));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam ss_i4_rep_411.GSR = "ENABLED";
    FD1P3IX dutyout_m1_i0_i9 (.D(n1258[9]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i9.GSR = "DISABLED";
    CCU2D add_179_15 (.A0(Out0[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18421), 
          .COUT(n18422), .S0(n1145[13]), .S1(n1145[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_15.INIT0 = 16'h5aaa;
    defparam add_179_15.INIT1 = 16'h5aaa;
    defparam add_179_15.INJECT1_0 = "NO";
    defparam add_179_15.INJECT1_1 = "NO";
    FD1P3IX dutyout_m1_i0_i8 (.D(n1258[8]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i7 (.D(n1258[7]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i7.GSR = "DISABLED";
    CCU2D add_15801_3 (.A0(speed_set_m3[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18673), .COUT(n18674));
    defparam add_15801_3.INIT0 = 16'hf555;
    defparam add_15801_3.INIT1 = 16'hf555;
    defparam add_15801_3.INJECT1_0 = "NO";
    defparam add_15801_3.INJECT1_1 = "NO";
    FD1P3IX dutyout_m1_i0_i6 (.D(n1258[6]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i6.GSR = "DISABLED";
    PFUMX addIn2_28__I_29_i13 (.BLUT(n618[12]), .ALUT(addIn2_28__N_1337[12]), 
          .C0(n20447), .Z(addIn2_28__N_1207[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    FD1P3IX dutyout_m1_i0_i5 (.D(n1258[5]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i4 (.D(n2152[4]), .SP(clk_N_683_enable_392), .CD(n12639), 
            .CK(clk_N_683), .Q(PWMdut_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i4.GSR = "DISABLED";
    CCU2D sub_16_rep_2_add_2_9 (.A0(subIn2[6]), .B0(n16636), .C0(n27[6]), 
          .D0(n2244[6]), .A1(subIn2[7]), .B1(n16636), .C1(n27[7]), .D1(n2244[7]), 
          .CIN(n18493), .COUT(n18494), .S0(subOut_24__N_1135[6]), .S1(subOut_24__N_1135[7]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_9.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_9.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_9.INJECT1_1 = "NO";
    LUT4 mux_137_i22_3_lut_4_lut_4_lut (.A(n21554), .B(n588[21]), .C(intgOut3[21]), 
         .D(n21552), .Z(n618[21])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i22_3_lut_4_lut_4_lut.init = 16'hccd8;
    CCU2D sub_16_rep_2_add_2_7 (.A0(subIn2[4]), .B0(n16636), .C0(n27[4]), 
          .D0(n2244[4]), .A1(subIn2[5]), .B1(n16636), .C1(n27[5]), .D1(n2244[5]), 
          .CIN(n18492), .COUT(n18493), .S0(subOut_24__N_1135[4]), .S1(subOut_24__N_1135[5]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_7.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_7.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_7.INJECT1_1 = "NO";
    FD1P3IX dutyout_m1_i0_i3 (.D(n1258[3]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i3.GSR = "DISABLED";
    PFUMX addIn2_28__I_29_i14 (.BLUT(n618[13]), .ALUT(addIn2_28__N_1337[13]), 
          .C0(n20447), .Z(addIn2_28__N_1207[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    FD1P3IX dutyout_m1_i0_i2 (.D(n2152[2]), .SP(clk_N_683_enable_392), .CD(n12639), 
            .CK(clk_N_683), .Q(PWMdut_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i2.GSR = "DISABLED";
    LUT4 mux_137_i23_3_lut_4_lut_4_lut (.A(n21554), .B(n588[22]), .C(intgOut3[22]), 
         .D(n21552), .Z(n618[22])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i23_3_lut_4_lut_4_lut.init = 16'hccd8;
    FD1P3IX dutyout_m1_i0_i1 (.D(n2152[1]), .SP(clk_N_683_enable_392), .CD(n12639), 
            .CK(clk_N_683), .Q(PWMdut_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m1_i0_i1.GSR = "DISABLED";
    PFUMX addIn2_28__I_29_i15 (.BLUT(n618[14]), .ALUT(addIn2_28__N_1337[14]), 
          .C0(n20447), .Z(addIn2_28__N_1207[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_137_i24_3_lut_4_lut_4_lut (.A(n21554), .B(n588[23]), .C(intgOut3[23]), 
         .D(n21552), .Z(n618[23])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i24_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX addIn2_28__I_29_i16 (.BLUT(n618[15]), .ALUT(addIn2_28__N_1337[15]), 
          .C0(n20447), .Z(addIn2_28__N_1207[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_137_i25_3_lut_4_lut_4_lut (.A(n21554), .B(n588[24]), .C(intgOut3[24]), 
         .D(n21552), .Z(n618[24])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i25_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX addIn2_28__I_29_i17 (.BLUT(n618[16]), .ALUT(addIn2_28__N_1337[16]), 
          .C0(n20447), .Z(addIn2_28__N_1207[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    LUT4 mux_137_i26_3_lut_4_lut_4_lut (.A(n21554), .B(n588[25]), .C(intgOut3[25]), 
         .D(n21552), .Z(n618[25])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i26_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX addIn2_28__I_29_i1 (.BLUT(n618[0]), .ALUT(addIn2_28__N_1337[0]), 
          .C0(n20447), .Z(addIn2_28__N_1207[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;
    CCU2D add_15801_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[0]), .B1(speed_set_m3[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18673));
    defparam add_15801_1.INIT0 = 16'hF000;
    defparam add_15801_1.INIT1 = 16'ha666;
    defparam add_15801_1.INJECT1_0 = "NO";
    defparam add_15801_1.INJECT1_1 = "NO";
    LUT4 mux_137_i27_3_lut_4_lut_4_lut (.A(n21554), .B(n588[26]), .C(intgOut3[26]), 
         .D(n21552), .Z(n618[26])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i27_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX mux_1801_i4 (.BLUT(n3690[3]), .ALUT(subIn2_24__N_1114[3]), .C0(n20179), 
          .Z(subIn2[3]));
    LUT4 mux_137_i28_3_lut_4_lut_4_lut (.A(n21554), .B(n588[27]), .C(intgOut3[27]), 
         .D(n21552), .Z(n618[27])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i28_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_137_i29_3_lut_4_lut_4_lut (.A(n21554), .B(n588[28]), .C(intgOut3[28]), 
         .D(n21552), .Z(n618[28])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_137_i29_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX mux_1801_i8 (.BLUT(n3690[7]), .ALUT(subIn2_24__N_1114[7]), .C0(n20179), 
          .Z(subIn2[7]));
    LUT4 i1_3_lut_4_lut_adj_76 (.A(n22208), .B(n920), .C(addOut[23]), 
         .D(n3635), .Z(intgOut0_28__N_735[23])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_76.init = 16'h1110;
    PFUMX mux_1801_i9 (.BLUT(n3690[8]), .ALUT(subIn2_24__N_1114[8]), .C0(n20179), 
          .Z(subIn2[8]));
    CCU2D add_179_13 (.A0(Out0[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18420), 
          .COUT(n18421), .S0(n1145[11]), .S1(n1145[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_13.INIT0 = 16'h5aaa;
    defparam add_179_13.INIT1 = 16'h5aaa;
    defparam add_179_13.INJECT1_0 = "NO";
    defparam add_179_13.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_77 (.A(n22208), .B(n920), .C(addOut[24]), 
         .D(n3635), .Z(intgOut0_28__N_735[24])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_77.init = 16'h1110;
    PFUMX mux_1801_i10 (.BLUT(n3690[9]), .ALUT(subIn2_24__N_1114[9]), .C0(n20179), 
          .Z(subIn2[9]));
    LUT4 i7_4_lut_adj_78 (.A(Out3[3]), .B(n14_adj_1837), .C(n10_adj_1838), 
         .D(Out3[4]), .Z(n18859)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam i7_4_lut_adj_78.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_79 (.A(n22208), .B(n920), .C(addOut[25]), 
         .D(n3635), .Z(intgOut0_28__N_735[25])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_79.init = 16'h1110;
    LUT4 i1_3_lut_4_lut_adj_80 (.A(n22208), .B(n920), .C(addOut[26]), 
         .D(n3635), .Z(intgOut0_28__N_735[26])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_80.init = 16'h1110;
    PFUMX mux_1801_i13 (.BLUT(n3690[12]), .ALUT(subIn2_24__N_1114[12]), 
          .C0(n20179), .Z(subIn2[12]));
    LUT4 i1_4_lut_adj_81 (.A(n21599), .B(n19740), .C(n22208), .D(n21583), 
         .Z(clk_N_683_enable_73)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_81.init = 16'hc4c0;
    LUT4 i1_3_lut_4_lut_adj_82 (.A(n22208), .B(n920), .C(addOut[27]), 
         .D(n3635), .Z(intgOut0_28__N_735[27])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_82.init = 16'h1110;
    LUT4 i1_3_lut_4_lut_adj_83 (.A(n22208), .B(n920), .C(addOut[28]), 
         .D(n3635), .Z(intgOut0_28__N_735[28])) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_83.init = 16'h1110;
    LUT4 mux_198_i4_3_lut_4_lut_3_lut (.A(n30_adj_1839), .B(n1145[15]), 
         .C(n2152[3]), .Z(n1258[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(326[25:42])
    defparam mux_198_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_198_i8_3_lut_4_lut_3_lut (.A(n30_adj_1839), .B(n1145[15]), 
         .C(n2152[7]), .Z(n1258[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(326[25:42])
    defparam mux_198_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    PFUMX mux_1801_i2 (.BLUT(subIn2_24__N_1301[1]), .ALUT(subIn2_24__N_1114[1]), 
          .C0(n20183), .Z(subIn2[1]));
    LUT4 mux_198_i10_3_lut_4_lut_3_lut (.A(n30_adj_1839), .B(n1145[15]), 
         .C(n2152[9]), .Z(n1258[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(326[25:42])
    defparam mux_198_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_198_i9_3_lut_4_lut_3_lut (.A(n30_adj_1839), .B(n1145[15]), 
         .C(n2152[8]), .Z(n1258[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(326[25:42])
    defparam mux_198_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_198_i7_3_lut_4_lut_3_lut (.A(n30_adj_1839), .B(n1145[15]), 
         .C(n2152[6]), .Z(n1258[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(326[25:42])
    defparam mux_198_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    CCU2D add_179_11 (.A0(Out0[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18419), 
          .COUT(n18420), .S0(n1145[9]), .S1(n1145[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_11.INIT0 = 16'h5aaa;
    defparam add_179_11.INIT1 = 16'h5aaa;
    defparam add_179_11.INJECT1_0 = "NO";
    defparam add_179_11.INJECT1_1 = "NO";
    PFUMX mux_1801_i3 (.BLUT(subIn2_24__N_1301[2]), .ALUT(subIn2_24__N_1114[2]), 
          .C0(n20183), .Z(subIn2[2]));
    LUT4 i1_2_lut_adj_84 (.A(ss[1]), .B(ss[2]), .Z(n19779)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_adj_84.init = 16'hbbbb;
    LUT4 mux_198_i6_3_lut_4_lut_3_lut (.A(n30_adj_1839), .B(n1145[15]), 
         .C(n2152[5]), .Z(n1258[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(326[25:42])
    defparam mux_198_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    PFUMX mux_1801_i5 (.BLUT(subIn2_24__N_1301[4]), .ALUT(subIn2_24__N_1114[4]), 
          .C0(n20183), .Z(subIn2[4]));
    CCU2D sub_16_rep_2_add_2_5 (.A0(subIn2[2]), .B0(n16636), .C0(n27[2]), 
          .D0(n2244[2]), .A1(subIn2[3]), .B1(n16636), .C1(n27[3]), .D1(n2244[3]), 
          .CIN(n18491), .COUT(n18492), .S0(subOut_24__N_1135[2]), .S1(subOut_24__N_1135[3]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_5.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_5.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_5.INJECT1_1 = "NO";
    PFUMX mux_1801_i6 (.BLUT(subIn2_24__N_1301[5]), .ALUT(subIn2_24__N_1114[5]), 
          .C0(n20183), .Z(subIn2[5]));
    CCU2D add_179_9 (.A0(Out0[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18418), 
          .COUT(n18419), .S0(n1145[7]), .S1(n1145[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_9.INIT0 = 16'h5aaa;
    defparam add_179_9.INIT1 = 16'h5aaa;
    defparam add_179_9.INJECT1_0 = "NO";
    defparam add_179_9.INJECT1_1 = "NO";
    LUT4 mux_138_i26_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[25]), 
         .D(intgOut2[25]), .Z(n648[25])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i26_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i10_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[9]), 
         .D(intgOut2[9]), .Z(n648[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i10_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15802_21 (.A0(speed_set_m1[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18672), .S1(n35));
    defparam add_15802_21.INIT0 = 16'h5555;
    defparam add_15802_21.INIT1 = 16'h0000;
    defparam add_15802_21.INJECT1_0 = "NO";
    defparam add_15802_21.INJECT1_1 = "NO";
    CCU2D add_15802_19 (.A0(speed_set_m1[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18671), .COUT(n18672));
    defparam add_15802_19.INIT0 = 16'hf555;
    defparam add_15802_19.INIT1 = 16'hf555;
    defparam add_15802_19.INJECT1_0 = "NO";
    defparam add_15802_19.INJECT1_1 = "NO";
    LUT4 mux_138_i9_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[8]), 
         .D(intgOut2[8]), .Z(n648[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i9_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i8_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[7]), 
         .D(intgOut2[7]), .Z(n648[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i29_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[28]), 
         .D(intgOut2[28]), .Z(n648[28])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i29_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i20_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[19]), 
         .D(intgOut2[19]), .Z(n648[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i20_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i21_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[20]), 
         .D(intgOut2[20]), .Z(n648[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i13_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[12]), 
         .D(intgOut2[12]), .Z(n648[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i11_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[10]), 
         .D(intgOut2[10]), .Z(n648[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i28_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[27]), 
         .D(intgOut2[27]), .Z(n648[27])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i28_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i27_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[26]), 
         .D(intgOut2[26]), .Z(n648[26])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i27_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i12_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[11]), 
         .D(intgOut2[11]), .Z(n648[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i12_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i22_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[21]), 
         .D(intgOut2[21]), .Z(n648[21])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i22_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i14_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[13]), 
         .D(intgOut2[13]), .Z(n648[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i14_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_179_7 (.A0(Out0[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18417), 
          .COUT(n18418), .S0(n1145[5]), .S1(n1145[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_7.INIT0 = 16'h5aaa;
    defparam add_179_7.INIT1 = 16'h5aaa;
    defparam add_179_7.INJECT1_0 = "NO";
    defparam add_179_7.INJECT1_1 = "NO";
    LUT4 mux_138_i2_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[1]), 
         .D(intgOut2[1]), .Z(n648[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i2_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15802_17 (.A0(speed_set_m1[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18670), .COUT(n18671));
    defparam add_15802_17.INIT0 = 16'hf555;
    defparam add_15802_17.INIT1 = 16'hf555;
    defparam add_15802_17.INJECT1_0 = "NO";
    defparam add_15802_17.INJECT1_1 = "NO";
    PFUMX mux_1801_i7 (.BLUT(subIn2_24__N_1301[6]), .ALUT(subIn2_24__N_1114[6]), 
          .C0(n20183), .Z(subIn2[6]));
    LUT4 mux_138_i23_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[22]), 
         .D(intgOut2[22]), .Z(n648[22])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i23_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i24_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[23]), 
         .D(intgOut2[23]), .Z(n648[23])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i24_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_179_5 (.A0(Out0[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18416), 
          .COUT(n18417), .S0(n1145[3]), .S1(n1145[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_5.INIT0 = 16'h5aaa;
    defparam add_179_5.INIT1 = 16'h5aaa;
    defparam add_179_5.INJECT1_0 = "NO";
    defparam add_179_5.INJECT1_1 = "NO";
    CCU2D sub_16_rep_2_add_2_3 (.A0(subIn2[0]), .B0(n16636), .C0(n27[0]), 
          .D0(n2244[0]), .A1(subIn2[1]), .B1(n16636), .C1(n27[1]), .D1(n2244[1]), 
          .CIN(n18490), .COUT(n18491), .S0(subOut_24__N_1135[0]), .S1(subOut_24__N_1135[1]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_3.INIT0 = 16'hb874;
    defparam sub_16_rep_2_add_2_3.INIT1 = 16'hb874;
    defparam sub_16_rep_2_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_3.INJECT1_1 = "NO";
    CCU2D add_179_3 (.A0(Out0[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18415), 
          .COUT(n18416), .S0(n1145[1]), .S1(n1145[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_3.INIT0 = 16'h5aaa;
    defparam add_179_3.INIT1 = 16'h5aaa;
    defparam add_179_3.INJECT1_0 = "NO";
    defparam add_179_3.INJECT1_1 = "NO";
    LUT4 mux_138_i15_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[14]), 
         .D(intgOut2[14]), .Z(n648[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 i2_3_lut_4_lut_adj_85 (.A(n15941), .B(n49), .C(n57), .D(n21490), 
         .Z(n16541)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(138[23] 139[51])
    defparam i2_3_lut_4_lut_adj_85.init = 16'hfff4;
    LUT4 mux_138_i16_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[15]), 
         .D(intgOut2[15]), .Z(n648[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_3_lut_4_lut_adj_86 (.A(n15941), .B(n49), .C(n16648), 
         .D(n21490), .Z(n2436)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(138[23] 139[51])
    defparam i1_2_lut_3_lut_4_lut_adj_86.init = 16'hf040;
    LUT4 i17063_2_lut (.A(ss[2]), .B(ss[1]), .Z(n19897)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17063_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_4_lut_adj_87 (.A(n21522), .B(n56), .C(n21486), .D(n21491), 
         .Z(n19788)) /* synthesis lut_function=(A (C+(D))+!A (B)) */ ;
    defparam i1_4_lut_4_lut_adj_87.init = 16'heee4;
    LUT4 mux_138_i25_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[24]), 
         .D(intgOut2[24]), .Z(n648[24])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i6_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[5]), 
         .D(intgOut2[5]), .Z(n648[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i7_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[6]), 
         .D(intgOut2[6]), .Z(n648[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i19_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[18]), 
         .D(intgOut2[18]), .Z(n648[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i19_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15802_15 (.A0(speed_set_m1[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18669), .COUT(n18670));
    defparam add_15802_15.INIT0 = 16'hf555;
    defparam add_15802_15.INIT1 = 16'hf555;
    defparam add_15802_15.INJECT1_0 = "NO";
    defparam add_15802_15.INJECT1_1 = "NO";
    LUT4 mux_138_i18_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[17]), 
         .D(intgOut2[17]), .Z(n648[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i18_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i17_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[16]), 
         .D(intgOut2[16]), .Z(n648[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i17_3_lut_4_lut.init = 16'hfe10;
    CCU2D sub_16_rep_2_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n19732), .B1(n21484), .C1(GND_net), .D1(GND_net), 
          .COUT(n18490));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_2_add_2_1.INIT0 = 16'hF000;
    defparam sub_16_rep_2_add_2_1.INIT1 = 16'h7777;
    defparam sub_16_rep_2_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_2_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_138_i3_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[2]), 
         .D(intgOut2[2]), .Z(n648[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i3_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_179_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[13]), .B1(n18864), .C1(n18865), .D1(Out0[28]), .COUT(n18415), 
          .S1(n1145[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(314[17:21])
    defparam add_179_1.INIT0 = 16'hF000;
    defparam add_179_1.INIT1 = 16'h56aa;
    defparam add_179_1.INJECT1_0 = "NO";
    defparam add_179_1.INJECT1_1 = "NO";
    LUT4 mux_138_i4_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[3]), 
         .D(intgOut2[3]), .Z(n648[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i5_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[4]), 
         .D(intgOut2[4]), .Z(n648[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i5_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i1_3_lut_4_lut (.A(n21552), .B(n21550), .C(intgOut1[0]), 
         .D(intgOut2[0]), .Z(n648[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(169[9:16])
    defparam mux_138_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_4_lut (.A(n22208), .B(n21607), .C(ss[3]), .D(ss[0]), 
         .Z(multIn2[6])) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h1400;
    LUT4 i17857_2_lut_rep_311_3_lut_3_lut_4_lut (.A(n22199), .B(n22196), 
         .C(n21584), .D(n21552), .Z(n21520)) /* synthesis lut_function=(!((B+!(C+!(D)))+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(165[9:16])
    defparam i17857_2_lut_rep_311_3_lut_3_lut_4_lut.init = 16'h2022;
    CCU2D add_15802_13 (.A0(speed_set_m1[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18668), .COUT(n18669));
    defparam add_15802_13.INIT0 = 16'hf555;
    defparam add_15802_13.INIT1 = 16'hf555;
    defparam add_15802_13.INJECT1_0 = "NO";
    defparam add_15802_13.INJECT1_1 = "NO";
    CCU2D add_15802_11 (.A0(speed_set_m1[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18667), .COUT(n18668));
    defparam add_15802_11.INIT0 = 16'hf555;
    defparam add_15802_11.INIT1 = 16'hf555;
    defparam add_15802_11.INJECT1_0 = "NO";
    defparam add_15802_11.INJECT1_1 = "NO";
    CCU2D add_15802_9 (.A0(speed_set_m1[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18666), .COUT(n18667));
    defparam add_15802_9.INIT0 = 16'hf555;
    defparam add_15802_9.INIT1 = 16'hf555;
    defparam add_15802_9.INJECT1_0 = "NO";
    defparam add_15802_9.INJECT1_1 = "NO";
    LUT4 i17867_2_lut_4_lut (.A(n22196), .B(n21584), .C(ss[2]), .D(n20579), 
         .Z(n20447)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(165[9:16])
    defparam i17867_2_lut_4_lut.init = 16'hff04;
    LUT4 i17855_2_lut_3_lut_4_lut (.A(n22196), .B(n21571), .C(n4138), 
         .D(ss[2]), .Z(n20183)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i17855_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i1_2_lut_rep_291_3_lut_4_lut_4_lut_4_lut (.A(n22199), .B(n21578), 
         .C(n21553), .D(n21552), .Z(n21500)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+!(D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(174[9:17])
    defparam i1_2_lut_rep_291_3_lut_4_lut_4_lut_4_lut.init = 16'h5051;
    LUT4 i13755_2_lut (.A(addOut[0]), .B(n22208), .Z(backOut1_28__N_1445[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13755_2_lut.init = 16'h2222;
    CCU2D add_1179_23 (.A0(n5177), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18414), 
          .S0(n2244[21]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_23.INIT0 = 16'hf555;
    defparam add_1179_23.INIT1 = 16'h0000;
    defparam add_1179_23.INJECT1_0 = "NO";
    defparam add_1179_23.INJECT1_1 = "NO";
    PFUMX mux_1801_i11 (.BLUT(subIn2_24__N_1301[10]), .ALUT(subIn2_24__N_1114[10]), 
          .C0(n20183), .Z(subIn2[10]));
    LUT4 i17844_2_lut_rep_276_2_lut (.A(n49), .B(n15941), .Z(n21485)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i17844_2_lut_rep_276_2_lut.init = 16'h1111;
    LUT4 mux_1244_i18_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[17]), 
         .C(speed_set_m3[17]), .D(n15941), .Z(n2484[17])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i18_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1244_i21_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[20]), 
         .C(speed_set_m3[20]), .D(n15941), .Z(n2484[20])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i21_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1244_i20_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[19]), 
         .C(speed_set_m3[19]), .D(n15941), .Z(n2484[19])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i20_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i1_4_lut_4_lut_4_lut_4_lut_3_lut_4_lut_4_lut (.A(n49), .B(n21484), 
         .C(n19788), .D(n15941), .Z(n19732)) /* synthesis lut_function=(A ((C)+!B)+!A ((C (D))+!B)) */ ;
    defparam i1_4_lut_4_lut_4_lut_4_lut_3_lut_4_lut_4_lut.init = 16'hf3b3;
    CCU2D add_15802_7 (.A0(speed_set_m1[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18665), .COUT(n18666));
    defparam add_15802_7.INIT0 = 16'hf555;
    defparam add_15802_7.INIT1 = 16'hf555;
    defparam add_15802_7.INJECT1_0 = "NO";
    defparam add_15802_7.INJECT1_1 = "NO";
    LUT4 i2_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n21485), .B(n21489), .C(n19788), 
         .D(n21487), .Z(n16636)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0040;
    CCU2D add_15802_5 (.A0(speed_set_m1[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18664), .COUT(n18665));
    defparam add_15802_5.INIT0 = 16'hf555;
    defparam add_15802_5.INIT1 = 16'hf555;
    defparam add_15802_5.INJECT1_0 = "NO";
    defparam add_15802_5.INJECT1_1 = "NO";
    CCU2D add_15802_3 (.A0(speed_set_m1[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18663), .COUT(n18664));
    defparam add_15802_3.INIT0 = 16'hf555;
    defparam add_15802_3.INIT1 = 16'hf555;
    defparam add_15802_3.INJECT1_0 = "NO";
    defparam add_15802_3.INJECT1_1 = "NO";
    CCU2D add_1179_21 (.A0(n5175), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5177), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18413), 
          .COUT(n18414), .S0(n2244[19]), .S1(n2244[20]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(126[13] 142[6])
    defparam add_1179_21.INIT0 = 16'hf555;
    defparam add_1179_21.INIT1 = 16'hf555;
    defparam add_1179_21.INJECT1_0 = "NO";
    defparam add_1179_21.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_88 (.A(ss[1]), .B(n19740), .C(n22208), .D(n19668), 
         .Z(clk_N_683_enable_325)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_88.init = 16'hc4c0;
    CCU2D add_15802_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[0]), .B1(speed_set_m1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18663));
    defparam add_15802_1.INIT0 = 16'hF000;
    defparam add_15802_1.INIT1 = 16'ha666;
    defparam add_15802_1.INJECT1_0 = "NO";
    defparam add_15802_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_89 (.A(ss[1]), .B(n19740), .C(n22208), .D(n19668), 
         .Z(clk_N_683_enable_353)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_89.init = 16'hc8c0;
    LUT4 mux_1244_i1_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[0]), .C(speed_set_m3[0]), 
         .D(n15941), .Z(n2484[0])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i1_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i13963_2_lut (.A(addOut[21]), .B(n22208), .Z(backOut1_28__N_1445[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13963_2_lut.init = 16'h2222;
    PFUMX mux_1801_i12 (.BLUT(subIn2_24__N_1301[11]), .ALUT(subIn2_24__N_1114[11]), 
          .C0(n20183), .Z(subIn2[11]));
    LUT4 i13962_2_lut (.A(addOut[20]), .B(n22208), .Z(backOut1_28__N_1445[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13962_2_lut.init = 16'h2222;
    CCU2D add_15810_21 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18593), .S1(n42));
    defparam add_15810_21.INIT0 = 16'h5555;
    defparam add_15810_21.INIT1 = 16'h0000;
    defparam add_15810_21.INJECT1_0 = "NO";
    defparam add_15810_21.INJECT1_1 = "NO";
    CCU2D add_15810_19 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18592), .COUT(n18593));
    defparam add_15810_19.INIT0 = 16'hf555;
    defparam add_15810_19.INIT1 = 16'hf555;
    defparam add_15810_19.INJECT1_0 = "NO";
    defparam add_15810_19.INJECT1_1 = "NO";
    CCU2D add_15810_17 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18591), .COUT(n18592));
    defparam add_15810_17.INIT0 = 16'hf555;
    defparam add_15810_17.INIT1 = 16'hf555;
    defparam add_15810_17.INJECT1_0 = "NO";
    defparam add_15810_17.INJECT1_1 = "NO";
    CCU2D add_15810_15 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18590), .COUT(n18591));
    defparam add_15810_15.INIT0 = 16'hf555;
    defparam add_15810_15.INIT1 = 16'hf555;
    defparam add_15810_15.INJECT1_0 = "NO";
    defparam add_15810_15.INJECT1_1 = "NO";
    CCU2D add_15810_13 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18589), .COUT(n18590));
    defparam add_15810_13.INIT0 = 16'hf555;
    defparam add_15810_13.INIT1 = 16'hf555;
    defparam add_15810_13.INJECT1_0 = "NO";
    defparam add_15810_13.INJECT1_1 = "NO";
    LUT4 i13953_2_lut (.A(addOut[19]), .B(n22208), .Z(backOut0_28__N_1416[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13953_2_lut.init = 16'h2222;
    LUT4 i13952_2_lut (.A(addOut[18]), .B(n22208), .Z(backOut0_28__N_1416[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13952_2_lut.init = 16'h2222;
    PFUMX mux_1801_i14 (.BLUT(subIn2_24__N_1301[13]), .ALUT(subIn2_24__N_1114[13]), 
          .C0(n20183), .Z(subIn2[13]));
    LUT4 i13951_2_lut (.A(addOut[17]), .B(n22208), .Z(backOut0_28__N_1416[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13951_2_lut.init = 16'h2222;
    LUT4 i13950_2_lut (.A(addOut[16]), .B(n22208), .Z(backOut0_28__N_1416[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13950_2_lut.init = 16'h2222;
    LUT4 i13949_2_lut (.A(addOut[15]), .B(n22208), .Z(backOut0_28__N_1416[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13949_2_lut.init = 16'h2222;
    LUT4 mux_1244_i19_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[18]), 
         .C(speed_set_m3[18]), .D(n15941), .Z(n2484[18])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i19_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i10230_3_lut_4_lut (.A(n1145[15]), .B(n30_adj_1839), .C(n18815), 
         .D(clk_N_683_enable_392), .Z(n12639)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(326[7:42])
    defparam i10230_3_lut_4_lut.init = 16'hf700;
    CCU2D add_15810_11 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18588), .COUT(n18589));
    defparam add_15810_11.INIT0 = 16'hf555;
    defparam add_15810_11.INIT1 = 16'hf555;
    defparam add_15810_11.INJECT1_0 = "NO";
    defparam add_15810_11.INJECT1_1 = "NO";
    CCU2D add_15810_9 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18587), .COUT(n18588));
    defparam add_15810_9.INIT0 = 16'hf555;
    defparam add_15810_9.INIT1 = 16'hf555;
    defparam add_15810_9.INJECT1_0 = "NO";
    defparam add_15810_9.INJECT1_1 = "NO";
    LUT4 i5_4_lut_adj_90 (.A(n9_adj_1840), .B(n7_adj_1841), .C(n1187[10]), 
         .D(n1187[13]), .Z(n30)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_90.init = 16'h8000;
    CCU2D add_15810_7 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18586), .COUT(n18587));
    defparam add_15810_7.INIT0 = 16'hf555;
    defparam add_15810_7.INIT1 = 16'hf555;
    defparam add_15810_7.INJECT1_0 = "NO";
    defparam add_15810_7.INJECT1_1 = "NO";
    LUT4 i3_2_lut_adj_91 (.A(n1187[14]), .B(n1187[12]), .Z(n9_adj_1840)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_91.init = 16'h8888;
    CCU2D add_15810_5 (.A0(speed_set_m2[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18585), .COUT(n18586));
    defparam add_15810_5.INIT0 = 16'hf555;
    defparam add_15810_5.INIT1 = 16'hf555;
    defparam add_15810_5.INJECT1_0 = "NO";
    defparam add_15810_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_92 (.A(n1187[11]), .B(n1187[9]), .C(n10_adj_1842), 
         .D(n1187[7]), .Z(n7_adj_1841)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_92.init = 16'haaa8;
    LUT4 i4_4_lut_adj_93 (.A(n1187[6]), .B(n8_adj_1843), .C(n1187[4]), 
         .D(n4_adj_1844), .Z(n10_adj_1842)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_93.init = 16'hfeee;
    LUT4 i2_2_lut_adj_94 (.A(n1187[5]), .B(n1187[8]), .Z(n8_adj_1843)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_94.init = 16'heeee;
    LUT4 i1_4_lut_adj_95 (.A(n1187[3]), .B(n1187[2]), .C(n1187[1]), .D(n1187[0]), 
         .Z(n4_adj_1844)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_95.init = 16'haaa8;
    LUT4 i13948_2_lut (.A(addOut[14]), .B(n22208), .Z(backOut0_28__N_1416[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13948_2_lut.init = 16'h2222;
    LUT4 i13947_2_lut (.A(addOut[13]), .B(n22208), .Z(backOut0_28__N_1416[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13947_2_lut.init = 16'h2222;
    LUT4 mux_1244_i17_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[16]), 
         .C(speed_set_m3[16]), .D(n15941), .Z(n2484[16])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i17_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX mux_1801_i15 (.BLUT(subIn2_24__N_1301[14]), .ALUT(subIn2_24__N_1114[14]), 
          .C0(n20183), .Z(subIn2[14]));
    LUT4 i13946_2_lut (.A(addOut[12]), .B(n22208), .Z(backOut0_28__N_1416[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13946_2_lut.init = 16'h2222;
    LUT4 i13961_2_lut (.A(addOut[11]), .B(n22208), .Z(backOut1_28__N_1445[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13961_2_lut.init = 16'h2222;
    LUT4 i13960_2_lut (.A(addOut[10]), .B(n22208), .Z(backOut1_28__N_1445[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13960_2_lut.init = 16'h2222;
    LUT4 i13959_2_lut (.A(addOut[9]), .B(n22208), .Z(backOut1_28__N_1445[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13959_2_lut.init = 16'h2222;
    LUT4 mux_1244_i16_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[15]), 
         .C(speed_set_m3[15]), .D(n15941), .Z(n2484[15])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i16_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i13956_2_lut (.A(addOut[28]), .B(n22208), .Z(backOut0_28__N_1416[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13956_2_lut.init = 16'h2222;
    LUT4 i13945_2_lut (.A(addOut[8]), .B(n22208), .Z(backOut0_28__N_1416[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13945_2_lut.init = 16'h2222;
    LUT4 i13944_2_lut (.A(addOut[7]), .B(n22208), .Z(backOut0_28__N_1416[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13944_2_lut.init = 16'h2222;
    LUT4 i13966_2_lut (.A(addOut[27]), .B(n22208), .Z(backOut1_28__N_1445[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13966_2_lut.init = 16'h2222;
    LUT4 mux_1244_i15_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[14]), 
         .C(speed_set_m3[14]), .D(n15941), .Z(n2484[14])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i15_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i13958_2_lut (.A(addOut[6]), .B(n22208), .Z(backOut1_28__N_1445[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13958_2_lut.init = 16'h2222;
    LUT4 i13957_2_lut (.A(addOut[5]), .B(n22208), .Z(backOut1_28__N_1445[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13957_2_lut.init = 16'h2222;
    LUT4 i13967_2_lut (.A(addOut[26]), .B(n22208), .Z(backOut2_28__N_1474[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13967_2_lut.init = 16'h2222;
    LUT4 mux_1244_i14_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[13]), 
         .C(speed_set_m3[13]), .D(n15941), .Z(n2484[13])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i14_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1244_i13_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[12]), 
         .C(speed_set_m3[12]), .D(n15941), .Z(n2484[12])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i13_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i13943_2_lut (.A(addOut[4]), .B(n22208), .Z(backOut0_28__N_1416[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13943_2_lut.init = 16'h2222;
    LUT4 i13942_2_lut (.A(addOut[3]), .B(n22208), .Z(backOut0_28__N_1416[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13942_2_lut.init = 16'h2222;
    LUT4 mux_1244_i12_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[11]), 
         .C(speed_set_m3[11]), .D(n15941), .Z(n2484[11])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i12_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1244_i11_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[10]), 
         .C(speed_set_m3[10]), .D(n15941), .Z(n2484[10])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i11_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1244_i10_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[9]), .C(speed_set_m3[9]), 
         .D(n15941), .Z(n2484[9])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i10_3_lut_4_lut_4_lut.init = 16'hccd8;
    CCU2D add_15810_3 (.A0(speed_set_m2[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18584), .COUT(n18585));
    defparam add_15810_3.INIT0 = 16'hf555;
    defparam add_15810_3.INIT1 = 16'hf555;
    defparam add_15810_3.INJECT1_0 = "NO";
    defparam add_15810_3.INJECT1_1 = "NO";
    LUT4 mux_1244_i9_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[8]), .C(speed_set_m3[8]), 
         .D(n15941), .Z(n2484[8])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i9_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1244_i8_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[7]), .C(speed_set_m3[7]), 
         .D(n15941), .Z(n2484[7])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i8_3_lut_4_lut_4_lut.init = 16'hccd8;
    CCU2D add_15810_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[0]), .B1(speed_set_m2[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18584));
    defparam add_15810_1.INIT0 = 16'hF000;
    defparam add_15810_1.INIT1 = 16'ha666;
    defparam add_15810_1.INJECT1_0 = "NO";
    defparam add_15810_1.INJECT1_1 = "NO";
    LUT4 mux_1244_i7_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[6]), .C(speed_set_m3[6]), 
         .D(n15941), .Z(n2484[6])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i7_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 i13941_2_lut (.A(addOut[2]), .B(n22208), .Z(backOut0_28__N_1416[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13941_2_lut.init = 16'h2222;
    LUT4 mux_1244_i6_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[5]), .C(speed_set_m3[5]), 
         .D(n15941), .Z(n2484[5])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i6_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1244_i5_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[4]), .C(speed_set_m3[4]), 
         .D(n15941), .Z(n2484[4])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i5_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX mux_1801_i16 (.BLUT(subIn2_24__N_1301[15]), .ALUT(subIn2_24__N_1114[15]), 
          .C0(n20183), .Z(subIn2[15]));
    CCU2D sub_16_rep_3_add_2_23 (.A0(n21486), .B0(n16648), .C0(n57), .D0(n5729), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18645), 
          .S0(n27[21]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_23.INIT0 = 16'h04ff;
    defparam sub_16_rep_3_add_2_23.INIT1 = 16'h0000;
    defparam sub_16_rep_3_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_23.INJECT1_1 = "NO";
    LUT4 mux_1244_i4_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[3]), .C(speed_set_m3[3]), 
         .D(n15941), .Z(n2484[3])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i4_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX mux_1801_i17 (.BLUT(subIn2_24__N_1301[16]), .ALUT(subIn2_24__N_1114[16]), 
          .C0(n20183), .Z(subIn2[16]));
    LUT4 mux_1244_i3_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[2]), .C(speed_set_m3[2]), 
         .D(n15941), .Z(n2484[2])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i3_3_lut_4_lut_4_lut.init = 16'hccd8;
    PFUMX mux_1801_i18 (.BLUT(subIn2_24__N_1301[17]), .ALUT(subIn2_24__N_1114[17]), 
          .C0(n20183), .Z(subIn2[17]));
    LUT4 mux_1244_i2_3_lut_4_lut_4_lut (.A(n49), .B(speed_set_m4[1]), .C(speed_set_m3[1]), 
         .D(n15941), .Z(n2484[1])) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mux_1244_i2_3_lut_4_lut_4_lut.init = 16'hccd8;
    LUT4 mux_1189_i1_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[0]), 
         .D(speed_set_m3[0]), .Z(n5045)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i1_3_lut_4_lut.init = 16'hfb40;
    CCU2D sub_16_rep_3_add_2_21 (.A0(n7), .B0(n16648), .C0(n16541), .D0(n5725), 
          .A1(n21486), .B1(n16648), .C1(n57), .D1(n5729), .CIN(n18644), 
          .COUT(n18645), .S0(n27[19]), .S1(n27[20]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_21.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_21.INIT1 = 16'h04ff;
    defparam sub_16_rep_3_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_21.INJECT1_1 = "NO";
    PFUMX mux_1801_i19 (.BLUT(subIn2_24__N_1301[18]), .ALUT(subIn2_24__N_1114[18]), 
          .C0(n20183), .Z(subIn2[18]));
    CCU2D add_191_17 (.A0(Out3[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18446), 
          .S0(n1208[15]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_17.INIT0 = 16'h5aaa;
    defparam add_191_17.INIT1 = 16'h0000;
    defparam add_191_17.INJECT1_0 = "NO";
    defparam add_191_17.INJECT1_1 = "NO";
    LUT4 i10232_3_lut_4_lut (.A(n1166[15]), .B(n30_adj_1833), .C(n18815), 
         .D(clk_N_683_enable_392), .Z(n12648)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(334[7:42])
    defparam i10232_3_lut_4_lut.init = 16'hf700;
    LUT4 i1_2_lut_rep_277_3_lut_4_lut (.A(n21499), .B(n42), .C(n49), .D(n15941), 
         .Z(n21486)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam i1_2_lut_rep_277_3_lut_4_lut.init = 16'h44f4;
    LUT4 mux_1189_i5_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[4]), 
         .D(speed_set_m3[4]), .Z(n5055)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i6_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[5]), 
         .D(speed_set_m3[5]), .Z(n5057)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1754_1_lut (.A(n42), .Z(subIn1_24__N_1300)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(137[34:50])
    defparam i1754_1_lut.init = 16'h5555;
    LUT4 i1755_1_lut (.A(n49), .Z(dirout_m3_N_1578)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(139[35:51])
    defparam i1755_1_lut.init = 16'h5555;
    CCU2D add_191_15 (.A0(Out3[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18445), 
          .COUT(n18446), .S0(n1208[13]), .S1(n1208[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_15.INIT0 = 16'h5aaa;
    defparam add_191_15.INIT1 = 16'h5aaa;
    defparam add_191_15.INJECT1_0 = "NO";
    defparam add_191_15.INJECT1_1 = "NO";
    LUT4 i1753_1_lut (.A(n35), .Z(subIn1_24__N_1113)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(135[34:50])
    defparam i1753_1_lut.init = 16'h5555;
    LUT4 i1756_1_lut (.A(n56), .Z(dirout_m4_N_1581)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(141[35:51])
    defparam i1756_1_lut.init = 16'h5555;
    LUT4 i13604_2_lut_rep_401 (.A(n22208), .B(ss[3]), .Z(n22196)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13604_2_lut_rep_401.init = 16'heeee;
    CCU2D add_191_13 (.A0(Out3[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18444), 
          .COUT(n18445), .S0(n1208[11]), .S1(n1208[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam add_191_13.INIT0 = 16'h5aaa;
    defparam add_191_13.INIT1 = 16'h5aaa;
    defparam add_191_13.INJECT1_0 = "NO";
    defparam add_191_13.INJECT1_1 = "NO";
    LUT4 mux_1189_i3_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[2]), 
         .D(speed_set_m3[2]), .Z(n5051)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i4_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[3]), 
         .D(speed_set_m3[3]), .Z(n5053)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i2_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[1]), 
         .D(speed_set_m3[1]), .Z(n5049)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i7_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[6]), 
         .D(speed_set_m3[6]), .Z(n5059)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i8_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[7]), 
         .D(speed_set_m3[7]), .Z(n5061)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i9_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[8]), 
         .D(speed_set_m3[8]), .Z(n5063)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i9_3_lut_4_lut.init = 16'hfb40;
    CCU2D sub_16_rep_3_add_2_19 (.A0(subIn2[17]), .B0(n16648), .C0(n16541), 
          .D0(n5721), .A1(subIn2[18]), .B1(n16648), .C1(n16541), .D1(n5723), 
          .CIN(n18643), .COUT(n18644), .S0(n27[17]), .S1(n27[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_19.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_19.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_19.INJECT1_1 = "NO";
    LUT4 mux_1189_i10_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[9]), 
         .D(speed_set_m3[9]), .Z(n5065)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i11_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[10]), 
         .D(speed_set_m3[10]), .Z(n5067)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i11_3_lut_4_lut.init = 16'hfb40;
    PFUMX mux_1801_i1 (.BLUT(subIn2_24__N_1301[0]), .ALUT(subIn2_24__N_1114[0]), 
          .C0(n20183), .Z(subIn2[0]));
    LUT4 mux_1188_i12_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m4[11]), .Z(n5111)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1189_i12_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[11]), 
         .D(speed_set_m3[11]), .Z(n5069)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i13_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[12]), 
         .D(speed_set_m3[12]), .Z(n5071)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i14_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[13]), 
         .D(speed_set_m3[13]), .Z(n5073)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i15_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[14]), 
         .D(speed_set_m3[14]), .Z(n5075)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i16_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[15]), 
         .D(speed_set_m3[15]), .Z(n5077)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i17_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[16]), 
         .D(speed_set_m3[16]), .Z(n5079)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i18_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[17]), 
         .D(speed_set_m3[17]), .Z(n5081)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i19_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[18]), 
         .D(speed_set_m3[18]), .Z(n5083)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i19_3_lut_4_lut.init = 16'hfb40;
    CCU2D sub_16_rep_3_add_2_17 (.A0(subIn2[15]), .B0(n16648), .C0(n16541), 
          .D0(n5717), .A1(subIn2[16]), .B1(n16648), .C1(n16541), .D1(n5719), 
          .CIN(n18642), .COUT(n18643), .S0(n27[15]), .S1(n27[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_17.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_17.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_15 (.A0(subIn2[13]), .B0(n16648), .C0(n16541), 
          .D0(n5713), .A1(subIn2[14]), .B1(n16648), .C1(n16541), .D1(n5715), 
          .CIN(n18641), .COUT(n18642), .S0(n27[13]), .S1(n27[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_15.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_15.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_15.INJECT1_1 = "NO";
    LUT4 mux_1189_i20_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[19]), 
         .D(speed_set_m3[19]), .Z(n5085)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1189_i21_3_lut_4_lut (.A(n21499), .B(n42), .C(speed_set_m2[20]), 
         .D(speed_set_m3[20]), .Z(n5087)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(136[23] 137[50])
    defparam mux_1189_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1188_i2_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m4[1]), .Z(n5091)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i2_3_lut_4_lut.init = 16'hf780;
    FD1P3IX dutyout_m4_i0_i9 (.D(n1390[9]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i8 (.D(n1390[8]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i7 (.D(n1390[7]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i6 (.D(n1390[6]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i5 (.D(n1390[5]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i4 (.D(n2188[4]), .SP(clk_N_683_enable_392), .CD(n12666), 
            .CK(clk_N_683), .Q(PWMdut_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i3 (.D(n1390[3]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i3.GSR = "DISABLED";
    CCU2D sub_16_rep_3_add_2_13 (.A0(subIn2[11]), .B0(n16648), .C0(n16541), 
          .D0(n5709), .A1(subIn2[12]), .B1(n16648), .C1(n16541), .D1(n5711), 
          .CIN(n18640), .COUT(n18641), .S0(n27[11]), .S1(n27[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_13.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_13.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_13.INJECT1_1 = "NO";
    FD1P3IX dutyout_m4_i0_i2 (.D(n2188[2]), .SP(clk_N_683_enable_392), .CD(n12666), 
            .CK(clk_N_683), .Q(PWMdut_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i1 (.D(n2188[1]), .SP(clk_N_683_enable_392), .CD(n12666), 
            .CK(clk_N_683), .Q(PWMdut_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i9 (.D(n1346[9]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i8 (.D(n1346[8]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i7 (.D(n1346[7]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i6 (.D(n1346[6]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i5 (.D(n1346[5]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i4 (.D(n2176[4]), .SP(clk_N_683_enable_392), .CD(n12655), 
            .CK(clk_N_683), .Q(PWMdut_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i3 (.D(n1346[3]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i2 (.D(n2176[2]), .SP(clk_N_683_enable_392), .CD(n12655), 
            .CK(clk_N_683), .Q(PWMdut_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i1 (.D(n2176[1]), .SP(clk_N_683_enable_392), .CD(n12655), 
            .CK(clk_N_683), .Q(PWMdut_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m3_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i9 (.D(n1302[9]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i8 (.D(n1302[8]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i7 (.D(n1302[7]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i6 (.D(n1302[6]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i5 (.D(n1302[5]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i5.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_adj_96 (.A(ss[1]), .B(n21583), .C(ss[3]), .D(n22208), 
         .Z(n19725)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut_adj_96.init = 16'h0080;
    FD1P3IX dutyout_m2_i0_i4 (.D(n2164[4]), .SP(clk_N_683_enable_392), .CD(n12648), 
            .CK(clk_N_683), .Q(PWMdut_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i3 (.D(n1302[3]), .SP(clk_N_683_enable_392), .CD(n12641), 
            .CK(clk_N_683), .Q(PWMdut_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i2 (.D(n2164[2]), .SP(clk_N_683_enable_392), .CD(n12648), 
            .CK(clk_N_683), .Q(PWMdut_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m2_i0_i2.GSR = "DISABLED";
    LUT4 mux_1188_i6_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m4[5]), .Z(n5099)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1188_i7_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m4[6]), .Z(n5101)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i13940_2_lut (.A(addOut[1]), .B(n22208), .Z(backOut0_28__N_1416[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13940_2_lut.init = 16'h2222;
    LUT4 mux_1188_i8_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m4[7]), .Z(n5103)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1188_i4_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m4[3]), .Z(n5095)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1188_i5_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m4[4]), .Z(n5097)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1188_i3_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m4[2]), .Z(n5093)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1188_i1_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m4[0]), .Z(n5047)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i1_3_lut_4_lut.init = 16'hf780;
    CCU2D sub_16_rep_3_add_2_11 (.A0(subIn2[9]), .B0(n16648), .C0(n16541), 
          .D0(n5705), .A1(subIn2[10]), .B1(n16648), .C1(n16541), .D1(n5707), 
          .CIN(n18639), .COUT(n18640), .S0(n27[9]), .S1(n27[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_11.INIT0 = 16'ha655;
    defparam sub_16_rep_3_add_2_11.INIT1 = 16'ha655;
    defparam sub_16_rep_3_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_11.INJECT1_1 = "NO";
    LUT4 mux_1188_i9_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m4[8]), .Z(n5105)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i6_4_lut_adj_97 (.A(Out3[11]), .B(Out3[7]), .C(Out3[2]), .D(Out3[10]), 
         .Z(n14_adj_1837)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam i6_4_lut_adj_97.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_98 (.A(n21608), .B(n21607), .C(n22203), 
         .D(n22208), .Z(n19740)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_3_lut_4_lut_adj_98.init = 16'he0f0;
    LUT4 mux_1188_i10_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m4[9]), .Z(n5107)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_2_lut_adj_99 (.A(Out3[9]), .B(Out3[1]), .Z(n10_adj_1838)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam i2_2_lut_adj_99.init = 16'heeee;
    LUT4 i4_4_lut_adj_100 (.A(Out3[5]), .B(Out3[6]), .C(Out3[0]), .D(n6_adj_1845), 
         .Z(n18860)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam i4_4_lut_adj_100.init = 16'hfffe;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n21608), .B(n21607), .C(n19897), .D(n22208), 
         .Z(clk_N_683_enable_129)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B !((D)+!C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_4_lut_4_lut_4_lut.init = 16'hee50;
    LUT4 i1_4_lut_4_lut_4_lut_adj_101 (.A(n21608), .B(n21607), .C(n19779), 
         .D(n22208), .Z(clk_N_683_enable_101)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_4_lut_4_lut_4_lut_adj_101.init = 16'hee05;
    LUT4 i1_2_lut_adj_102 (.A(Out3[8]), .B(Out3[12]), .Z(n6_adj_1845)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(317[17:21])
    defparam i1_2_lut_adj_102.init = 16'heeee;
    LUT4 i13965_2_lut (.A(addOut[25]), .B(n22208), .Z(backOut1_28__N_1445[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13965_2_lut.init = 16'h2222;
    LUT4 i1838_2_lut_rep_362 (.A(ss[0]), .B(ss[1]), .Z(n21571)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1838_2_lut_rep_362.init = 16'h6666;
    LUT4 i1_2_lut_rep_321_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n22199), 
         .D(n22196), .Z(n21530)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_321_3_lut_4_lut.init = 16'h0006;
    LUT4 mux_1188_i13_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m4[12]), .Z(n5113)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i13955_2_lut (.A(addOut[24]), .B(n22208), .Z(backOut0_28__N_1416[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13955_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_335_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n22199), 
         .D(n22196), .Z(n21544)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_rep_335_3_lut_4_lut.init = 16'h0060;
    LUT4 i13954_2_lut (.A(addOut[23]), .B(n22208), .Z(backOut0_28__N_1416[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13954_2_lut.init = 16'h2222;
    LUT4 i1814_1_lut_rep_363 (.A(ss[0]), .Z(n21572)) /* synthesis lut_function=(!(A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1814_1_lut_rep_363.init = 16'h5555;
    LUT4 equal_114_i6_2_lut_rep_343_2_lut (.A(ss[0]), .B(ss[1]), .Z(n21552)) /* synthesis lut_function=((B)+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam equal_114_i6_2_lut_rep_343_2_lut.init = 16'hdddd;
    LUT4 equal_114_i9_2_lut_rep_315_3_lut_4_lut_4_lut (.A(ss[0]), .B(ss[2]), 
         .C(n21578), .D(ss[1]), .Z(n21524)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam equal_114_i9_2_lut_rep_315_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i17979_2_lut_rep_301_2_lut_3_lut_4_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21578), .D(n22199), .Z(n21510)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i17979_2_lut_rep_301_2_lut_3_lut_4_lut_4_lut.init = 16'h0002;
    LUT4 ss_4__I_0_319_i9_2_lut_rep_334_3_lut_4_lut_4_lut (.A(ss[0]), .B(ss[2]), 
         .C(n22196), .D(ss[1]), .Z(n21543)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam ss_4__I_0_319_i9_2_lut_rep_334_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_4_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(n21607), .D(n22208), 
         .Z(n4147)) /* synthesis lut_function=(!(A+(B (C+(D))+!B ((D)+!C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h0014;
    LUT4 i1_4_lut_4_lut_then_4_lut (.A(ss[1]), .B(ss[2]), .C(ss[3]), .D(ss[0]), 
         .Z(n21610)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_4_lut_then_4_lut.init = 16'hfffe;
    LUT4 ss_4__I_0_317_i9_2_lut_rep_320_3_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21578), .D(ss[2]), .Z(n21529)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(192[19:27])
    defparam ss_4__I_0_317_i9_2_lut_rep_320_3_lut_4_lut.init = 16'hfffb;
    LUT4 i5_4_lut_adj_103 (.A(n9_adj_1846), .B(n7_adj_1847), .C(n1166[10]), 
         .D(n1166[13]), .Z(n30_adj_1833)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_103.init = 16'h8000;
    LUT4 mux_1188_i14_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m4[13]), .Z(n5115)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i17982_2_lut_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21578), 
         .D(n22199), .Z(n15859)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(192[19:27])
    defparam i17982_2_lut_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 ss_4__I_0_314_i6_2_lut_rep_368 (.A(ss[0]), .B(ss[1]), .Z(n21577)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(165[9:16])
    defparam ss_4__I_0_314_i6_2_lut_rep_368.init = 16'heeee;
    LUT4 i1_3_lut_rep_300_4_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21554), 
         .D(n21550), .Z(n21509)) /* synthesis lut_function=(A+(B (C)+!B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(172[20:27])
    defparam i1_3_lut_rep_300_4_lut_4_lut.init = 16'hfbea;
    LUT4 i3_2_lut_adj_104 (.A(n1166[14]), .B(n1166[12]), .Z(n9_adj_1846)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_104.init = 16'h8888;
    LUT4 i1_2_lut_rep_369 (.A(n22208), .B(ss[3]), .Z(n21578)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(174[9:17])
    defparam i1_2_lut_rep_369.init = 16'hbbbb;
    CCU2D add_15798_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18717), 
          .S0(n920));
    defparam add_15798_cout.INIT0 = 16'h0000;
    defparam add_15798_cout.INIT1 = 16'h0000;
    defparam add_15798_cout.INJECT1_0 = "NO";
    defparam add_15798_cout.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_340_3_lut (.A(n22208), .B(ss[3]), .C(n22199), .Z(n21549)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(174[9:17])
    defparam i1_2_lut_rep_340_3_lut.init = 16'hbfbf;
    CCU2D add_15798_22 (.A0(addOut[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18716), .COUT(n18717));
    defparam add_15798_22.INIT0 = 16'h5555;
    defparam add_15798_22.INIT1 = 16'hf555;
    defparam add_15798_22.INJECT1_0 = "NO";
    defparam add_15798_22.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_345_3_lut (.A(n22208), .B(ss[3]), .C(ss[2]), .Z(n21554)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(174[9:17])
    defparam i1_2_lut_rep_345_3_lut.init = 16'hfbfb;
    LUT4 equal_110_i9_2_lut_rep_319_3_lut_4_lut (.A(n22208), .B(ss[3]), 
         .C(n21584), .D(n22199), .Z(n21528)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(174[9:17])
    defparam equal_110_i9_2_lut_rep_319_3_lut_4_lut.init = 16'hffbf;
    LUT4 i1_4_lut_adj_105 (.A(n1166[11]), .B(n1166[9]), .C(n10_adj_1848), 
         .D(n1166[7]), .Z(n7_adj_1847)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_105.init = 16'haaa8;
    LUT4 mux_1188_i15_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m4[14]), .Z(n5117)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1188_i16_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m4[15]), .Z(n5119)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i16_3_lut_4_lut.init = 16'hf780;
    CCU2D add_15798_20 (.A0(addOut[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18715), .COUT(n18716));
    defparam add_15798_20.INIT0 = 16'h5555;
    defparam add_15798_20.INIT1 = 16'h5555;
    defparam add_15798_20.INJECT1_0 = "NO";
    defparam add_15798_20.INJECT1_1 = "NO";
    CCU2D add_15798_18 (.A0(addOut[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18714), .COUT(n18715));
    defparam add_15798_18.INIT0 = 16'h5555;
    defparam add_15798_18.INIT1 = 16'h5555;
    defparam add_15798_18.INJECT1_0 = "NO";
    defparam add_15798_18.INJECT1_1 = "NO";
    CCU2D add_15798_16 (.A0(addOut[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18713), .COUT(n18714));
    defparam add_15798_16.INIT0 = 16'h5555;
    defparam add_15798_16.INIT1 = 16'h5555;
    defparam add_15798_16.INJECT1_0 = "NO";
    defparam add_15798_16.INJECT1_1 = "NO";
    CCU2D add_15798_14 (.A0(addOut[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18712), .COUT(n18713));
    defparam add_15798_14.INIT0 = 16'h5aaa;
    defparam add_15798_14.INIT1 = 16'h5555;
    defparam add_15798_14.INJECT1_0 = "NO";
    defparam add_15798_14.INJECT1_1 = "NO";
    LUT4 mux_1188_i17_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m4[16]), .Z(n5121)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i4_4_lut_adj_106 (.A(n1166[6]), .B(n8_adj_1849), .C(n1166[4]), 
         .D(n4_adj_1850), .Z(n10_adj_1848)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_106.init = 16'hfeee;
    LUT4 mux_1188_i18_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m4[17]), .Z(n5123)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i2_2_lut_adj_107 (.A(n1166[5]), .B(n1166[8]), .Z(n8_adj_1849)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_107.init = 16'heeee;
    FD1P3IX dutyout_m4_i0_i0 (.D(n2188[0]), .SP(clk_N_683_enable_392), .CD(n12666), 
            .CK(clk_N_683), .Q(PWMdut_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=297, LSE_RLINE=297 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam dutyout_m4_i0_i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_108 (.A(n1166[3]), .B(n1166[2]), .C(n1166[1]), .D(n1166[0]), 
         .Z(n4_adj_1850)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_108.init = 16'haaa8;
    LUT4 ss_4__I_0_321_i9_2_lut_rep_317_3_lut_4_lut (.A(n22208), .B(ss[3]), 
         .C(n21584), .D(n22199), .Z(n21526)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam ss_4__I_0_321_i9_2_lut_rep_317_3_lut_4_lut.init = 16'hefff;
    LUT4 mux_1188_i19_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m4[18]), .Z(n5125)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 i5_4_lut_adj_109 (.A(n9_adj_1851), .B(n7_adj_1852), .C(n1145[10]), 
         .D(n1145[13]), .Z(n30_adj_1839)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_109.init = 16'h8000;
    LUT4 i3_2_lut_adj_110 (.A(n1145[14]), .B(n1145[12]), .Z(n9_adj_1851)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_110.init = 16'h8888;
    LUT4 i1_2_lut_rep_341_3_lut (.A(n22208), .B(ss[3]), .C(ss[2]), .Z(n21550)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_341_3_lut.init = 16'hefef;
    LUT4 i17994_3_lut_rep_342_4_lut (.A(n22208), .B(ss[3]), .C(n22199), 
         .D(n21584), .Z(n21551)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i17994_3_lut_rep_342_4_lut.init = 16'h0100;
    LUT4 mux_1188_i20_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m4[19]), .Z(n5127)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(n22208), .B(ss[3]), .C(ss[1]), 
         .D(ss[0]), .Z(n21553)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'h0110;
    LUT4 i1_4_lut_adj_111 (.A(n1145[11]), .B(n1145[9]), .C(n10_adj_1853), 
         .D(n1145[7]), .Z(n7_adj_1852)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_111.init = 16'haaa8;
    LUT4 i4_4_lut_adj_112 (.A(n1145[6]), .B(n8_adj_1854), .C(n1145[4]), 
         .D(n4_adj_1855), .Z(n10_adj_1853)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_112.init = 16'hfeee;
    LUT4 i2_2_lut_adj_113 (.A(n1145[5]), .B(n1145[8]), .Z(n8_adj_1854)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_113.init = 16'heeee;
    LUT4 mux_1188_i21_3_lut_4_lut (.A(n21500), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m4[20]), .Z(n5129)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(134[23] 135[50])
    defparam mux_1188_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_114 (.A(n1145[3]), .B(n1145[2]), .C(n1145[1]), .D(n1145[0]), 
         .Z(n4_adj_1855)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_114.init = 16'haaa8;
    FD1S3IX ss_i2_rep_402 (.D(n14), .CK(clk_N_683), .CD(ss[4]), .Q(n22199));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(204[2] 392[9])
    defparam ss_i2_rep_402.GSR = "ENABLED";
    LUT4 i13964_2_lut (.A(addOut[22]), .B(n22208), .Z(backOut1_28__N_1445[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(235[3] 390[12])
    defparam i13964_2_lut.init = 16'h2222;
    FD1S3AX addOut_2063__i1 (.D(n121[1]), .CK(clk_N_683), .Q(addOut[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i1.GSR = "ENABLED";
    PFUMX i18140 (.BLUT(n21612), .ALUT(n21613), .C0(ss[0]), .Z(n4132));
    FD1S3AX addOut_2063__i2 (.D(n121[2]), .CK(clk_N_683), .Q(addOut[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i2.GSR = "ENABLED";
    FD1S3AX addOut_2063__i3 (.D(n121[3]), .CK(clk_N_683), .Q(addOut[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i3.GSR = "ENABLED";
    FD1S3AX addOut_2063__i4 (.D(n121[4]), .CK(clk_N_683), .Q(addOut[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i4.GSR = "ENABLED";
    FD1S3AX addOut_2063__i5 (.D(n121[5]), .CK(clk_N_683), .Q(addOut[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i5.GSR = "ENABLED";
    FD1S3AX addOut_2063__i6 (.D(n121[6]), .CK(clk_N_683), .Q(addOut[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i6.GSR = "ENABLED";
    FD1S3AX addOut_2063__i7 (.D(n121[7]), .CK(clk_N_683), .Q(addOut[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i7.GSR = "ENABLED";
    FD1S3AX addOut_2063__i8 (.D(n121[8]), .CK(clk_N_683), .Q(addOut[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i8.GSR = "ENABLED";
    FD1S3AX addOut_2063__i9 (.D(n121[9]), .CK(clk_N_683), .Q(addOut[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i9.GSR = "ENABLED";
    FD1S3AX addOut_2063__i10 (.D(n121[10]), .CK(clk_N_683), .Q(addOut[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i10.GSR = "ENABLED";
    FD1S3AX addOut_2063__i11 (.D(n121[11]), .CK(clk_N_683), .Q(addOut[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i11.GSR = "ENABLED";
    FD1S3AX addOut_2063__i12 (.D(n121[12]), .CK(clk_N_683), .Q(addOut[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i12.GSR = "ENABLED";
    FD1S3AX addOut_2063__i13 (.D(n121[13]), .CK(clk_N_683), .Q(addOut[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i13.GSR = "ENABLED";
    FD1S3AX addOut_2063__i14 (.D(n121[14]), .CK(clk_N_683), .Q(addOut[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i14.GSR = "ENABLED";
    FD1S3AX addOut_2063__i15 (.D(n121[15]), .CK(clk_N_683), .Q(addOut[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i15.GSR = "ENABLED";
    FD1S3AX addOut_2063__i16 (.D(n121[16]), .CK(clk_N_683), .Q(addOut[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i16.GSR = "ENABLED";
    FD1S3AX addOut_2063__i17 (.D(n121[17]), .CK(clk_N_683), .Q(addOut[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i17.GSR = "ENABLED";
    FD1S3AX addOut_2063__i18 (.D(n121[18]), .CK(clk_N_683), .Q(addOut[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i18.GSR = "ENABLED";
    FD1S3AX addOut_2063__i19 (.D(n121[19]), .CK(clk_N_683), .Q(addOut[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i19.GSR = "ENABLED";
    FD1S3AX addOut_2063__i20 (.D(n121[20]), .CK(clk_N_683), .Q(addOut[20])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i20.GSR = "ENABLED";
    FD1S3AX addOut_2063__i21 (.D(n121[21]), .CK(clk_N_683), .Q(addOut[21])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i21.GSR = "ENABLED";
    FD1S3AX addOut_2063__i22 (.D(n121[22]), .CK(clk_N_683), .Q(addOut[22])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i22.GSR = "ENABLED";
    FD1S3AX addOut_2063__i23 (.D(n121[23]), .CK(clk_N_683), .Q(addOut[23])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i23.GSR = "ENABLED";
    FD1S3AX addOut_2063__i24 (.D(n121[24]), .CK(clk_N_683), .Q(addOut[24])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i24.GSR = "ENABLED";
    FD1S3AX addOut_2063__i25 (.D(n121[25]), .CK(clk_N_683), .Q(addOut[25])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i25.GSR = "ENABLED";
    FD1S3AX addOut_2063__i26 (.D(n121[26]), .CK(clk_N_683), .Q(addOut[26])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i26.GSR = "ENABLED";
    FD1S3AX addOut_2063__i27 (.D(n121[27]), .CK(clk_N_683), .Q(addOut[27])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i27.GSR = "ENABLED";
    FD1S3AX addOut_2063__i28 (.D(n121[28]), .CK(clk_N_683), .Q(addOut[28])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pid.vhd(230[13:19])
    defparam addOut_2063__i28.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR
//

module PWMGENERATOR (PWM_m4, pwm_clk, free_m4, clkout_c_enable_176, 
            hallsense_m4, n21587, enable_m4, n3223, n21589, n3187, 
            PWMdut_m4, GND_net);
    output PWM_m4;
    input pwm_clk;
    output free_m4;
    input clkout_c_enable_176;
    input [2:0]hallsense_m4;
    output n21587;
    input enable_m4;
    output n3223;
    output n21589;
    output n3187;
    input [9:0]PWMdut_m4;
    input GND_net;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_1805, free_N_1817, n18521;
    wire [9:0]cnt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(41[10:13])
    
    wire n3687, n18520, n7, n18519, n18518, n9, n10, n18517, 
        n12550;
    wire [9:0]n45;
    
    wire n10_adj_1824, n10959, n18541, n18540, n18539, n18538, n18537, 
        n14, n10_adj_1825, n19977, n6, n19997;
    
    FD1S3AX PWM_20 (.D(PWM_N_1805), .CK(pwm_clk), .Q(PWM_m4)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=338, LSE_RLINE=338 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1817), .SP(clkout_c_enable_176), .CK(pwm_clk), 
            .Q(free_m4));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i1721_3_lut_rep_378 (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .Z(n21587)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1721_3_lut_rep_378.init = 16'h1414;
    LUT4 i17951_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .D(enable_m4), .Z(n3223)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17951_2_lut_4_lut.init = 16'hebff;
    LUT4 i1691_3_lut_rep_380 (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .Z(n21589)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i1691_3_lut_rep_380.init = 16'h1414;
    LUT4 i17948_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .D(enable_m4), .Z(n3187)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(52[2] 76[9])
    defparam i17948_2_lut_4_lut.init = 16'hebff;
    CCU2D sub_1795_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m4[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18521), .S1(n3687));
    defparam sub_1795_add_2_11.INIT0 = 16'h5999;
    defparam sub_1795_add_2_11.INIT1 = 16'h0000;
    defparam sub_1795_add_2_11.INJECT1_0 = "NO";
    defparam sub_1795_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1795_add_2_9 (.A0(PWMdut_m4[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m4[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18520), 
          .COUT(n18521));
    defparam sub_1795_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1795_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1795_add_2_9.INJECT1_0 = "NO";
    defparam sub_1795_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1795_add_2_7 (.A0(PWMdut_m4[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m4[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18519), 
          .COUT(n18520));
    defparam sub_1795_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1795_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1795_add_2_7.INJECT1_0 = "NO";
    defparam sub_1795_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1795_add_2_5 (.A0(PWMdut_m4[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m4[4]), .C1(n9), .D1(n10), .CIN(n18518), 
          .COUT(n18519));
    defparam sub_1795_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1795_add_2_5.INIT1 = 16'h5999;
    defparam sub_1795_add_2_5.INJECT1_0 = "NO";
    defparam sub_1795_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1795_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m4[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m4[2]), .C1(n9), .D1(n10), .CIN(n18517), 
          .COUT(n18518));
    defparam sub_1795_add_2_3.INIT0 = 16'h5999;
    defparam sub_1795_add_2_3.INIT1 = 16'h5999;
    defparam sub_1795_add_2_3.INJECT1_0 = "NO";
    defparam sub_1795_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1795_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m4[0]), .C1(n9), .D1(n10), 
          .COUT(n18517));
    defparam sub_1795_add_2_1.INIT0 = 16'h0000;
    defparam sub_1795_add_2_1.INIT1 = 16'h5999;
    defparam sub_1795_add_2_1.INJECT1_0 = "NO";
    defparam sub_1795_add_2_1.INJECT1_1 = "NO";
    FD1S3IX cnt_2067__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n12550), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i1.GSR = "ENABLED";
    LUT4 i2_3_lut (.A(PWMdut_m4[5]), .B(PWMdut_m4[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_1824), .B(PWMdut_m4[9]), .C(PWMdut_m4[8]), 
         .D(PWMdut_m4[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2256_3_lut (.A(n10959), .B(PWMdut_m4[4]), .C(PWMdut_m4[3]), 
         .Z(n10_adj_1824)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2256_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D cnt_2067_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18541), .S0(n45[9]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2067_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18540), 
          .COUT(n18541), .S0(n45[7]), .S1(n45[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18539), 
          .COUT(n18540), .S0(n45[5]), .S1(n45[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18538), 
          .COUT(n18539), .S0(n45[3]), .S1(n45[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2067_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18537), 
          .COUT(n18538), .S0(n45[1]), .S1(n45[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2067_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2067_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_3.INJECT1_1 = "NO";
    LUT4 i1797_1_lut (.A(n3687), .Z(PWM_N_1805)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1797_1_lut.init = 16'h5555;
    CCU2D cnt_2067_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18537), .S1(n45[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2067_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2067_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2067_add_4_1.INJECT1_1 = "NO";
    LUT4 i17891_4_lut (.A(PWMdut_m4[5]), .B(n14), .C(n10_adj_1825), .D(PWMdut_m4[8]), 
         .Z(free_N_1817)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i17891_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m4[9]), .B(PWMdut_m4[3]), .C(PWMdut_m4[4]), 
         .D(n10959), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[7]), .Z(n10_adj_1825)) /* synthesis lut_function=(A+(B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_42 (.A(PWMdut_m4[2]), .B(PWMdut_m4[1]), .C(PWMdut_m4[0]), 
         .Z(n10959)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_42.init = 16'hfefe;
    LUT4 i17143_4_lut (.A(cnt[7]), .B(cnt[5]), .C(cnt[9]), .D(cnt[3]), 
         .Z(n19977)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17143_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(cnt[4]), .B(cnt[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i17163_3_lut (.A(cnt[6]), .B(n19977), .C(cnt[8]), .Z(n19997)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17163_3_lut.init = 16'h8080;
    LUT4 i17894_4_lut (.A(cnt[2]), .B(n19997), .C(cnt[1]), .D(n6), .Z(n12550)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(73[6:16])
    defparam i17894_4_lut.init = 16'h0004;
    FD1S3IX cnt_2067__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n12550), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i0.GSR = "ENABLED";
    FD1S3IX cnt_2067__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n12550), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i2.GSR = "ENABLED";
    FD1S3IX cnt_2067__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n12550), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i3.GSR = "ENABLED";
    FD1S3IX cnt_2067__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n12550), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i4.GSR = "ENABLED";
    FD1S3IX cnt_2067__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n12550), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i5.GSR = "ENABLED";
    FD1S3IX cnt_2067__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n12550), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i6.GSR = "ENABLED";
    FD1S3IX cnt_2067__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n12550), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i7.GSR = "ENABLED";
    FD1S3IX cnt_2067__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n12550), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i8.GSR = "ENABLED";
    FD1S3IX cnt_2067__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n12550), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/pwm_gen.vhd(72[9:12])
    defparam cnt_2067__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module HALL
//

module HALL (clk_1mhz, \speed_m4[0] , clkout_c_enable_176, hallsense_m4, 
            HALL_A_OUT_c_c, HALL_B_OUT_c_c, HALL_C_OUT_c_c, clkout_c_enable_164, 
            \speed_m4[1] , \speed_m4[2] , \speed_m4[3] , \speed_m4[4] , 
            \speed_m4[5] , \speed_m4[6] , \speed_m4[7] , \speed_m4[8] , 
            \speed_m4[9] , \speed_m4[10] , \speed_m4[11] , \speed_m4[12] , 
            \speed_m4[13] , \speed_m4[14] , \speed_m4[15] , \speed_m4[16] , 
            \speed_m4[17] , \speed_m4[18] , \speed_m4[19] , GND_net, 
            n22198);
    input clk_1mhz;
    output \speed_m4[0] ;
    input clkout_c_enable_176;
    output [2:0]hallsense_m4;
    input HALL_A_OUT_c_c;
    input HALL_B_OUT_c_c;
    input HALL_C_OUT_c_c;
    input clkout_c_enable_164;
    output \speed_m4[1] ;
    output \speed_m4[2] ;
    output \speed_m4[3] ;
    output \speed_m4[4] ;
    output \speed_m4[5] ;
    output \speed_m4[6] ;
    output \speed_m4[7] ;
    output \speed_m4[8] ;
    output \speed_m4[9] ;
    output \speed_m4[10] ;
    output \speed_m4[11] ;
    output \speed_m4[12] ;
    output \speed_m4[13] ;
    output \speed_m4[14] ;
    output \speed_m4[15] ;
    output \speed_m4[16] ;
    output \speed_m4[17] ;
    output \speed_m4[18] ;
    output \speed_m4[19] ;
    input GND_net;
    input n22198;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1mhz */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/toplevelfinal.vhd(86[9:17])
    wire [19:0]speedt;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_47, n4329;
    wire [19:0]n7;
    wire [6:0]stable_count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(62[10:22])
    
    wire stable_counting, n21492;
    wire [6:0]stable_counting_N_1759;
    wire [19:0]speedt_19__N_1678;
    
    wire hall3_old, hall3_lat, hall1_lat, hall2_lat, hall1_old, hall2_old, 
        n19645, n18842, stable_counting_N_1746, n21495, n21504, n21503, 
        n21518, n21542, n21519, n19877, n21541;
    wire [19:0]count;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(60[10:15])
    
    wire n5227, n21602, n21564, n21540, n21603, n13_adj_1818, n11_adj_1819, 
        n19096, n54, n17124, n19941, n20_adj_1820, n32, n19943, 
        n4, n19689, n17_adj_1821, n16_adj_1822, n12_adj_1823, n18486, 
        n18485, n18484, n18483, n18482, n18481, n18480, n18479, 
        n18478, n18477;
    
    FD1P3IX speedt__i0 (.D(n7[0]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i0.GSR = "ENABLED";
    FD1P3IX stable_count__i0 (.D(stable_counting_N_1759[0]), .SP(stable_counting), 
            .CD(n21492), .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1678[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall3_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall1_lat_57 (.D(HALL_A_OUT_c_c), .SP(clkout_c_enable_176), 
            .CK(clk_1mhz), .Q(hall1_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(HALL_B_OUT_c_c), .SP(clkout_c_enable_176), 
            .CK(clk_1mhz), .Q(hall2_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(HALL_C_OUT_c_c), .SP(clkout_c_enable_176), 
            .CK(clk_1mhz), .Q(hall3_lat));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_176), .CK(clk_1mhz), 
            .Q(hall1_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_164), .CK(clk_1mhz), 
            .Q(hall2_old));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 i2_3_lut_rep_286 (.A(n19645), .B(n18842), .C(stable_counting_N_1746), 
         .Z(n21495)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_286.init = 16'hfefe;
    LUT4 i2202_2_lut_rep_283_4_lut (.A(n19645), .B(n18842), .C(stable_counting_N_1746), 
         .D(stable_counting), .Z(n21492)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2202_2_lut_rep_283_4_lut.init = 16'h0100;
    LUT4 i3_3_lut_4_lut (.A(n21504), .B(n21503), .C(n21518), .D(n21542), 
         .Z(n18842)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[7:23])
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    LUT4 i13879_2_lut_4_lut (.A(stable_count[6]), .B(stable_count[5]), .C(n21519), 
         .D(stable_counting_N_1746), .Z(stable_counting_N_1759[6])) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (((D)+!C)+!B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13879_2_lut_4_lut.init = 16'h006a;
    LUT4 i17043_2_lut_3_lut_4_lut (.A(stable_count[5]), .B(n21519), .C(n21542), 
         .D(n21503), .Z(n19877)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i17043_2_lut_3_lut_4_lut.init = 16'hfff6;
    FD1P3IX speedt__i1 (.D(n7[1]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i1.GSR = "ENABLED";
    FD1P3IX speedt__i2 (.D(n7[2]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i2.GSR = "ENABLED";
    FD1P3IX speedt__i3 (.D(n7[3]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i3.GSR = "ENABLED";
    FD1P3IX speedt__i4 (.D(n7[4]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i4.GSR = "ENABLED";
    FD1P3IX speedt__i5 (.D(n7[5]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i5.GSR = "ENABLED";
    FD1P3IX speedt__i6 (.D(n7[6]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i6.GSR = "ENABLED";
    FD1P3IX speedt__i7 (.D(n7[7]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i7.GSR = "ENABLED";
    FD1P3IX speedt__i8 (.D(n7[8]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i8.GSR = "ENABLED";
    FD1P3IX speedt__i9 (.D(n7[9]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i9.GSR = "ENABLED";
    FD1P3IX speedt__i10 (.D(n7[10]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i10.GSR = "ENABLED";
    FD1P3IX speedt__i11 (.D(n7[11]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i11.GSR = "ENABLED";
    FD1P3IX speedt__i12 (.D(n7[12]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i12.GSR = "ENABLED";
    FD1P3IX speedt__i13 (.D(n7[13]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i13.GSR = "ENABLED";
    FD1P3IX speedt__i14 (.D(n7[14]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i14.GSR = "ENABLED";
    FD1P3IX speedt__i15 (.D(n7[15]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i15.GSR = "ENABLED";
    FD1P3IX speedt__i16 (.D(n7[16]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i16.GSR = "ENABLED";
    FD1P3IX speedt__i17 (.D(n7[17]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i17.GSR = "ENABLED";
    FD1P3IX speedt__i18 (.D(n7[18]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i18.GSR = "ENABLED";
    FD1P3IX speedt__i19 (.D(n7[19]), .SP(clk_1mhz_enable_47), .CD(n4329), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speedt__i19.GSR = "ENABLED";
    LUT4 i2496_3_lut_rep_294_4_lut (.A(stable_count[4]), .B(n21541), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n21503)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2496_3_lut_rep_294_4_lut.init = 16'h7f80;
    LUT4 i13878_2_lut_3_lut_4_lut (.A(stable_count[4]), .B(n21541), .C(stable_counting_N_1746), 
         .D(stable_count[5]), .Z(stable_counting_N_1759[5])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13878_2_lut_3_lut_4_lut.init = 16'h0708;
    FD1S3IX count__i1 (.D(n7[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n7[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n7[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n7[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n7[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n7[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n7[7]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n7[8]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n7[9]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n7[10]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(n7[11]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n7[12]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n7[13]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n7[14]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n7[15]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(n7[16]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(n7[17]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(n7[18]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(n7[19]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(stable_counting_N_1759[1]), .SP(stable_counting), 
            .CD(n21492), .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(stable_counting_N_1759[2]), .SP(stable_counting), 
            .CD(n21492), .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(stable_counting_N_1759[3]), .SP(stable_counting), 
            .CD(n21492), .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(stable_counting_N_1759[4]), .SP(stable_counting), 
            .CD(n21492), .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(stable_counting_N_1759[5]), .SP(stable_counting), 
            .CD(n21492), .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i6 (.D(stable_counting_N_1759[6]), .SP(stable_counting), 
            .CD(n21492), .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3AX speed__i2 (.D(speedt_19__N_1678[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1678[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1678[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1678[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1678[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1678[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1678[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1678[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1678[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1678[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1678[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1678[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1678[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1678[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1678[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1678[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1678[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1678[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1678[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i17884_4_lut (.A(stable_counting_N_1746), .B(stable_counting), 
         .C(n18842), .D(n19645), .Z(n5227)) /* synthesis lut_function=(A (B)+!A !((C+(D))+!B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(97[3] 113[10])
    defparam i17884_4_lut.init = 16'h888c;
    LUT4 i1_2_lut_rep_393 (.A(stable_count[0]), .B(stable_count[1]), .Z(n21602)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_2_lut_rep_393.init = 16'h8888;
    LUT4 i2470_2_lut_rep_355_3_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[2]), .Z(n21564)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i2470_2_lut_rep_355_3_lut.init = 16'h8080;
    LUT4 mux_28_i2_4_lut (.A(n7[1]), .B(speedt[1]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i2_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i3_4_lut (.A(n7[2]), .B(speedt[2]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i3_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i4_4_lut (.A(n7[3]), .B(speedt[3]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i4_4_lut.init = 16'hcaa0;
    LUT4 i13875_2_lut_3_lut_4_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_counting_N_1746), .D(stable_count[2]), .Z(stable_counting_N_1759[2])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i13875_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 mux_28_i5_4_lut (.A(n7[4]), .B(speedt[4]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i5_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i6_4_lut (.A(n7[5]), .B(speedt[5]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i6_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i7_4_lut (.A(n7[6]), .B(speedt[6]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i7_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i8_4_lut (.A(n7[7]), .B(speedt[7]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i8_4_lut.init = 16'hcaa0;
    LUT4 i2477_2_lut_rep_332_3_lut_4_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21541)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i2477_2_lut_rep_332_3_lut_4_lut.init = 16'h8000;
    LUT4 i2475_2_lut_rep_333_3_lut_4_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21542)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i2475_2_lut_rep_333_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2468_2_lut_rep_394 (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[2]), .Z(n21603)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i2468_2_lut_rep_394.init = 16'h7878;
    LUT4 stable_count_0__bdd_4_lut_4_lut (.A(stable_count[0]), .B(stable_count[1]), 
         .C(stable_count[2]), .D(stable_counting_N_1746), .Z(n19645)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_count_0__bdd_4_lut_4_lut.init = 16'h99fd;
    LUT4 mux_28_i9_4_lut (.A(n7[8]), .B(speedt[8]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i9_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i10_4_lut (.A(n7[9]), .B(speedt[9]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i10_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i11_4_lut (.A(n7[10]), .B(speedt[10]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i11_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i12_4_lut (.A(n7[11]), .B(speedt[11]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i12_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i13_4_lut (.A(n7[12]), .B(speedt[12]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i13_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i14_4_lut (.A(n7[13]), .B(speedt[13]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i14_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i15_4_lut (.A(n7[14]), .B(speedt[14]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i15_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i16_4_lut (.A(n7[15]), .B(speedt[15]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i16_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i17_4_lut (.A(n7[16]), .B(speedt[16]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i17_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i18_4_lut (.A(n7[17]), .B(speedt[17]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i18_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i19_4_lut (.A(n7[18]), .B(speedt[18]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i19_4_lut.init = 16'hcaa0;
    LUT4 mux_28_i20_4_lut (.A(n7[19]), .B(speedt[19]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i20_4_lut.init = 16'hcaa0;
    LUT4 i17888_3_lut (.A(n21540), .B(n21495), .C(stable_counting), .Z(clk_1mhz_enable_47)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(97[3] 113[10])
    defparam i17888_3_lut.init = 16'h7575;
    LUT4 i7_4_lut (.A(n13_adj_1818), .B(n11_adj_1819), .C(count[2]), .D(n19096), 
         .Z(n4329)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[5]), .B(n54), .C(stable_counting), .D(stable_counting_N_1746), 
         .Z(n13_adj_1818)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i5_4_lut.init = 16'h0080;
    LUT4 i1_4_lut (.A(clk_1mhz_enable_47), .B(n17124), .C(n19941), .D(n20_adj_1820), 
         .Z(n19096)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(62[10:22])
    defparam i1_4_lut.init = 16'h0800;
    LUT4 i17107_4_lut (.A(count[15]), .B(count[10]), .C(count[11]), .D(count[8]), 
         .Z(n19941)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17107_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(n32), .B(n19943), .C(count[0]), .D(count[13]), 
         .Z(n20_adj_1820)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i9_4_lut.init = 16'h0002;
    LUT4 i1_4_lut_adj_36 (.A(n19877), .B(stable_counting_N_1746), .C(n21603), 
         .D(n21518), .Z(n32)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i1_4_lut_adj_36.init = 16'hcccd;
    LUT4 i17109_4_lut (.A(count[6]), .B(stable_counting_N_1759[0]), .C(count[12]), 
         .D(count[7]), .Z(n19943)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17109_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_37 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_37.init = 16'h7bde;
    LUT4 i1_4_lut_rep_331 (.A(n54), .B(n19689), .C(count[2]), .D(count[5]), 
         .Z(n21540)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i1_4_lut_rep_331.init = 16'hdfff;
    LUT4 i13877_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21564), .C(stable_counting_N_1746), 
         .D(stable_count[4]), .Z(stable_counting_N_1759[4])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13877_2_lut_3_lut_4_lut.init = 16'h0708;
    LUT4 i2489_2_lut_rep_295_3_lut_4_lut (.A(stable_count[3]), .B(n21564), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21504)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2489_2_lut_rep_295_3_lut_4_lut.init = 16'h78f0;
    LUT4 i9_4_lut_adj_38 (.A(n17_adj_1821), .B(count[11]), .C(n16_adj_1822), 
         .D(n11_adj_1819), .Z(n19689)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i9_4_lut_adj_38.init = 16'hfeff;
    LUT4 i7_4_lut_adj_39 (.A(count[7]), .B(count[8]), .C(count[10]), .D(count[15]), 
         .Z(n17_adj_1821)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_39.init = 16'hfffe;
    LUT4 i6_4_lut (.A(count[13]), .B(count[12]), .C(count[6]), .D(count[0]), 
         .Z(n16_adj_1822)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[3]), .B(count[1]), .Z(n11_adj_1819)) /* synthesis lut_function=(A (B)) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_40 (.A(count[4]), .B(n12_adj_1823), .C(count[18]), 
         .D(count[9]), .Z(n54)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i6_4_lut_adj_40.init = 16'h8000;
    LUT4 i5_4_lut_adj_41 (.A(count[14]), .B(count[19]), .C(count[17]), 
         .D(count[16]), .Z(n12_adj_1823)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam i5_4_lut_adj_41.init = 16'h8000;
    LUT4 i24_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n17124)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(62[10:22])
    defparam i24_2_lut.init = 16'h6666;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18486), 
          .S0(n7[19]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18485), .COUT(n18486), .S0(n7[17]), .S1(n7[18]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18484), .COUT(n18485), .S0(n7[15]), .S1(n7[16]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    LUT4 mux_28_i1_4_lut (.A(n7[0]), .B(speedt[0]), .C(n21495), .D(n21540), 
         .Z(speedt_19__N_1678[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(105[4] 111[11])
    defparam mux_28_i1_4_lut.init = 16'hcaa0;
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18483), .COUT(n18484), .S0(n7[13]), .S1(n7[14]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18482), .COUT(n18483), .S0(n7[11]), .S1(n7[12]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18481), .COUT(n18482), .S0(n7[9]), .S1(n7[10]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18480), 
          .COUT(n18481), .S0(n7[7]), .S1(n7[8]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18479), 
          .COUT(n18480), .S0(n7[5]), .S1(n7[6]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18478), 
          .COUT(n18479), .S0(n7[3]), .S1(n7[4]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_354 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(stable_counting_N_1746)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_354.init = 16'hdede;
    LUT4 i17880_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .D(stable_count[0]), 
         .Z(stable_counting_N_1759[0])) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C+(D))))) */ ;
    defparam i17880_2_lut_4_lut.init = 16'h0021;
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18477), 
          .COUT(n18478), .S0(n7[1]), .S1(n7[2]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .D(n17124), 
         .Z(stable_counting_N_1759[1])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 i2482_2_lut_rep_309_3_lut_4_lut (.A(stable_count[2]), .B(n21602), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21518)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2482_2_lut_rep_309_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2484_2_lut_rep_310_3_lut_4_lut (.A(stable_count[2]), .B(n21602), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21519)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i2484_2_lut_rep_310_3_lut_4_lut.init = 16'h8000;
    LUT4 i13876_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21602), .C(stable_counting_N_1746), 
         .D(stable_count[3]), .Z(stable_counting_N_1759[3])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(99[21:33])
    defparam i13876_2_lut_3_lut_4_lut.init = 16'h0708;
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18477), 
          .S1(n7[0]));   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    FD1P3IX stable_counting_62 (.D(n22198), .SP(stable_counting_N_1746), 
            .CD(n5227), .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(n7[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_47), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // d:/wybedata/projects/roboteamtwente/electronics/lattice/motorcontroller/hallinput.vhd(75[2] 120[9])
    defparam count__i0.GSR = "ENABLED";
    
endmodule
