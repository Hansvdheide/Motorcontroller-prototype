// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.8.0.115.3
// Netlist written on Mon Jun 26 11:00:38 2017
//
// Verilog Description of module SPI_loopback_Top
//

module SPI_loopback_Top (CS, SCK, MOSI, MISO, HALL_A_OUT, HALL_B_OUT, 
            HALL_C_OUT, LED1, LED2, LED3, LED4, clkout, H_A_m1, 
            H_B_m1, H_C_m1, MA_m1, MB_m1, MC_m1, H_A_m2, H_B_m2, 
            H_C_m2, MA_m2, MB_m2, MC_m2, H_A_m3, H_B_m3, H_C_m3, 
            MA_m3, MB_m3, MC_m3, H_A_m4, H_B_m4, H_C_m4, MA_m4, 
            MB_m4, MC_m4);   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(24[8:24])
    input CS;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(27[2:4])
    input SCK;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(28[2:5])
    input MOSI;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(29[2:6])
    output MISO;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(30[2:6])
    output HALL_A_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(33[2:12])
    output HALL_B_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(34[2:12])
    output HALL_C_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(35[2:12])
    output LED1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(38[2:6])
    output LED2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(39[2:6])
    output LED3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(40[2:6])
    output LED4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(41[2:6])
    output clkout;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    input H_A_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(47[2:8])
    input H_B_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(48[2:8])
    input H_C_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(49[2:8])
    output [1:0]MA_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    output [1:0]MB_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    output [1:0]MC_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    input H_A_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(55[2:8])
    input H_B_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(56[2:8])
    input H_C_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(57[2:8])
    output [1:0]MA_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    output [1:0]MB_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    output [1:0]MC_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    input H_A_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(63[2:8])
    input H_B_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(64[2:8])
    input H_C_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(65[2:8])
    output [1:0]MA_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    output [1:0]MB_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    output [1:0]MC_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    input H_A_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(71[2:8])
    input H_B_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(72[2:8])
    input H_C_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(73[2:8])
    output [1:0]MA_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    output [1:0]MB_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    output [1:0]MC_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    wire clk_N_875 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    
    wire GND_net, VCC_net, CS_c, SCK_c, MOSI_c, HALL_A_OUT_c_c, 
        HALL_B_OUT_c_c, HALL_C_OUT_c_c, LED1_c, LED2_c, LED3_c, LED4_c, 
        MA_m1_c_1, MA_m1_c_0, MB_m1_c_1, MB_m1_c_0, MC_m1_c_1, MC_m1_c_0, 
        H_A_m2_c, H_B_m2_c, H_C_m2_c, MA_m2_c_1, MA_m2_c_0, MB_m2_c_1, 
        MB_m2_c_0, MC_m2_c_1, MC_m2_c_0, H_A_m3_c, H_B_m3_c, H_C_m3_c, 
        MA_m3_c_1, MA_m3_c_0, MB_m3_c_1, MB_m3_c_0, MC_m3_c_1, MC_m3_c_0, 
        H_A_m4_c, H_B_m4_c, H_C_m4_c, MA_m4_c_1, MA_m4_c_0, MB_m4_c_1, 
        MB_m4_c_0, MC_m4_c_1, MC_m4_c_0, rst, enable_m1, enable_m2, 
        enable_m3, enable_m4;
    wire [20:0]speed_set_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(99[9:21])
    wire [20:0]speed_set_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(100[9:21])
    wire [20:0]speed_set_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(101[9:21])
    wire [20:0]speed_set_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(102[9:21])
    wire [20:0]speed_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(104[9:17])
    wire [20:0]speed_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(105[9:17])
    wire [20:0]speed_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(106[9:17])
    wire [20:0]speed_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(107[9:17])
    wire [2:0]hallsense_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(110[9:21])
    wire [2:0]hallsense_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(111[9:21])
    wire [2:0]hallsense_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(112[9:21])
    wire [2:0]hallsense_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(113[9:21])
    
    wire PWM_m1, PWM_m2, PWM_m3, PWM_m4;
    wire [9:0]PWMdut_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(120[9:18])
    wire [9:0]PWMdut_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(121[9:18])
    wire [9:0]PWMdut_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(122[9:18])
    wire [9:0]PWMdut_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(123[9:18])
    
    wire dir_m1, dir_m2, dir_m3, dir_m4;
    wire [13:0]start_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(135[9:18])
    
    wire free_m1, free_m2, free_m3, free_m4;
    wire [20:0]speed_avg_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(144[9:21])
    wire [20:0]speed_avg_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(145[9:21])
    wire [20:0]speed_avg_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(146[9:21])
    wire [20:0]speed_avg_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(147[9:21])
    
    wire n3290, n3232, n3196, n3244, n3208, n3182, n3124, n19830, 
        n3088, n3136, n3100, n3074, n3016, n2980, n3028, n2992, 
        n2966, n2908, MISO_N_816, n4497, n4494, n4467, n4460, 
        n2884, n19843, n4498;
    wire [25:0]subOut_24__N_1369;
    
    wire n4499, n4500, n2872, n4490, n4487, n4484, n4481, n4471, 
        n4464, n4457, n4455, n18896, n18836, n6, n19826, n22430, 
        n2920, n4475, n4474, n4473, n4472, n4470, n4469, n4468, 
        n4466, n4465, n4463, n4462, n4461, n4459, n4458, n4456, 
        n4454, n4453, n18900, n4496, n4495, n4493, n4492, n4491, 
        n4489, n4488, n4486, n4485, n4483, n4482, n4480, n4479, 
        n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
        n72, n73, n74, n75, n18539, n18538, n18537, n18536, 
        n18535, n18534, n18533, n5172, n10424, n21649, clkout_c_enable_341, 
        clkout_c_enable_272, n22435, n19942, n21716, n21714, n21713, 
        n21712, n21710, n21709, clkout_c_enable_362, n21705, n21703, 
        n21702, n21700, n19845, n21696, n21695;
    
    VHI i2 (.Z(VCC_net));
    OSCH OSCInst0 (.STDBY(GND_net), .OSC(clkout_c)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCInst0.NOM_FREQ = "38.00";
    LUT4 m1_lut (.Z(n22430)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    FD1S3AX rst_12_rep_426 (.D(n21649), .CK(clkout_c), .Q(n22435));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12_rep_426.GSR = "DISABLED";
    OB MA_m2_pad_0 (.I(MA_m2_c_0), .O(MA_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    FD1P3AX start_cnt_2097__i0 (.D(n75), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i0.GSR = "DISABLED";
    OB HALL_B_OUT_pad (.I(HALL_B_OUT_c_c), .O(HALL_B_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(34[2:12])
    OB HALL_A_OUT_pad (.I(HALL_A_OUT_c_c), .O(HALL_A_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(33[2:12])
    OB MA_m2_pad_1 (.I(MA_m2_c_1), .O(MA_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    IB HALL_B_OUT_c_pad (.I(H_B_m1), .O(HALL_B_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(48[2:8])
    OBZ n5171_pad (.I(MISO_N_816), .T(n5172), .O(MISO));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    IB HALL_A_OUT_c_pad (.I(H_A_m1), .O(HALL_A_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(47[2:8])
    IB MOSI_pad (.I(MOSI), .O(MOSI_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(29[2:6])
    IB SCK_pad (.I(SCK), .O(SCK_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(28[2:5])
    IB CS_pad (.I(CS), .O(CS_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(27[2:4])
    OB MC_m4_pad_0 (.I(MC_m4_c_0), .O(MC_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    OB MC_m4_pad_1 (.I(MC_m4_c_1), .O(MC_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    OB MB_m4_pad_0 (.I(MB_m4_c_0), .O(MB_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    OB MB_m4_pad_1 (.I(MB_m4_c_1), .O(MB_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    OB MC_m1_pad_0 (.I(MC_m1_c_0), .O(MC_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    OB MC_m1_pad_1 (.I(MC_m1_c_1), .O(MC_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    OB MA_m4_pad_0 (.I(MA_m4_c_0), .O(MA_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_0 (.I(MB_m1_c_0), .O(MB_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    OB MA_m4_pad_1 (.I(MA_m4_c_1), .O(MA_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_1 (.I(MB_m1_c_1), .O(MB_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    OB MC_m3_pad_0 (.I(MC_m3_c_0), .O(MC_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    IB H_C_m4_pad (.I(H_C_m4), .O(H_C_m4_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(73[2:8])
    OB MA_m1_pad_0 (.I(MA_m1_c_0), .O(MA_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    OB MC_m3_pad_1 (.I(MC_m3_c_1), .O(MC_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    IB H_B_m4_pad (.I(H_B_m4), .O(H_B_m4_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(72[2:8])
    OB MA_m1_pad_1 (.I(MA_m1_c_1), .O(MA_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    OB MB_m3_pad_0 (.I(MB_m3_c_0), .O(MB_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    IB H_A_m4_pad (.I(H_A_m4), .O(H_A_m4_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(71[2:8])
    OB clkout_pad (.I(clkout_c), .O(clkout));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    OB MB_m3_pad_1 (.I(MB_m3_c_1), .O(MB_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    IB H_C_m3_pad (.I(H_C_m3), .O(H_C_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(65[2:8])
    OB LED4_pad (.I(LED4_c), .O(LED4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(41[2:6])
    OB MA_m3_pad_0 (.I(MA_m3_c_0), .O(MA_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    IB H_B_m3_pad (.I(H_B_m3), .O(H_B_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(64[2:8])
    OB LED3_pad (.I(LED3_c), .O(LED3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(40[2:6])
    OB MA_m3_pad_1 (.I(MA_m3_c_1), .O(MA_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    IB H_A_m3_pad (.I(H_A_m3), .O(H_A_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(63[2:8])
    OB LED2_pad (.I(LED2_c), .O(LED2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(39[2:6])
    OB MC_m2_pad_0 (.I(MC_m2_c_0), .O(MC_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    IB H_C_m2_pad (.I(H_C_m2), .O(H_C_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(57[2:8])
    OB LED1_pad (.I(LED1_c), .O(LED1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(38[2:6])
    OB MC_m2_pad_1 (.I(MC_m2_c_1), .O(MC_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    IB H_B_m2_pad (.I(H_B_m2), .O(H_B_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(56[2:8])
    OB HALL_C_OUT_pad (.I(HALL_C_OUT_c_c), .O(HALL_C_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(35[2:12])
    OB MB_m2_pad_0 (.I(MB_m2_c_0), .O(MB_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    IB H_A_m2_pad (.I(H_A_m2), .O(H_A_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(55[2:8])
    OB MB_m2_pad_1 (.I(MB_m2_c_1), .O(MB_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    IB HALL_C_OUT_c_pad (.I(H_C_m1), .O(HALL_C_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(49[2:8])
    LUT4 mux_2169_i1_3_lut (.A(n4475), .B(n4500), .C(n19942), .Z(subOut_24__N_1369[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i1_3_lut.init = 16'hacac;
    CCU2D start_cnt_2097_add_4_15 (.A0(start_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18539), .S0(n62));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_15.INIT0 = 16'hfaaa;
    defparam start_cnt_2097_add_4_15.INIT1 = 16'h0000;
    defparam start_cnt_2097_add_4_15.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_15.INJECT1_1 = "NO";
    CCU2D start_cnt_2097_add_4_13 (.A0(start_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18538), .COUT(n18539), .S0(n64), .S1(n63));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_13.INIT0 = 16'hfaaa;
    defparam start_cnt_2097_add_4_13.INIT1 = 16'hfaaa;
    defparam start_cnt_2097_add_4_13.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_13.INJECT1_1 = "NO";
    LUT4 i7927_2_lut (.A(n21649), .B(n62), .Z(n10424)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam i7927_2_lut.init = 16'heeee;
    CCU2D start_cnt_2097_add_4_11 (.A0(start_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18537), .COUT(n18538), .S0(n66), .S1(n65));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_11.INIT0 = 16'hfaaa;
    defparam start_cnt_2097_add_4_11.INIT1 = 16'hfaaa;
    defparam start_cnt_2097_add_4_11.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_11.INJECT1_1 = "NO";
    CCU2D start_cnt_2097_add_4_9 (.A0(start_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18536), .COUT(n18537), .S0(n68), .S1(n67));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_9.INIT0 = 16'hfaaa;
    defparam start_cnt_2097_add_4_9.INIT1 = 16'hfaaa;
    defparam start_cnt_2097_add_4_9.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_9.INJECT1_1 = "NO";
    CCU2D start_cnt_2097_add_4_7 (.A0(start_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18535), .COUT(n18536), .S0(n70), .S1(n69));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_7.INIT0 = 16'hfaaa;
    defparam start_cnt_2097_add_4_7.INIT1 = 16'hfaaa;
    defparam start_cnt_2097_add_4_7.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_7.INJECT1_1 = "NO";
    CCU2D start_cnt_2097_add_4_5 (.A0(start_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18534), .COUT(n18535), .S0(n72), .S1(n71));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_5.INIT0 = 16'hfaaa;
    defparam start_cnt_2097_add_4_5.INIT1 = 16'hfaaa;
    defparam start_cnt_2097_add_4_5.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_5.INJECT1_1 = "NO";
    CCU2D start_cnt_2097_add_4_3 (.A0(start_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18533), .COUT(n18534), .S0(n74), .S1(n73));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_3.INIT0 = 16'hfaaa;
    defparam start_cnt_2097_add_4_3.INIT1 = 16'hfaaa;
    defparam start_cnt_2097_add_4_3.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_3.INJECT1_1 = "NO";
    CCU2D start_cnt_2097_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18533), .S1(n75));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097_add_4_1.INIT0 = 16'hF000;
    defparam start_cnt_2097_add_4_1.INIT1 = 16'h0555;
    defparam start_cnt_2097_add_4_1.INJECT1_0 = "NO";
    defparam start_cnt_2097_add_4_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut (.A(n18900), .B(start_cnt[10]), .C(start_cnt[9]), .D(start_cnt[8]), 
         .Z(n18836)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_202 (.A(n18896), .B(n6), .C(start_cnt[6]), .D(start_cnt[4]), 
         .Z(n18900)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_202.init = 16'hfefc;
    LUT4 i3_4_lut_adj_203 (.A(start_cnt[0]), .B(start_cnt[3]), .C(start_cnt[2]), 
         .D(start_cnt[1]), .Z(n18896)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_203.init = 16'hfffe;
    LUT4 i2_2_lut (.A(start_cnt[7]), .B(start_cnt[5]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 mux_2169_i2_3_lut (.A(n4474), .B(n4499), .C(n19942), .Z(subOut_24__N_1369[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i2_3_lut.init = 16'hacac;
    LUT4 mux_2169_i3_3_lut (.A(n4473), .B(n4498), .C(n19942), .Z(subOut_24__N_1369[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i3_3_lut.init = 16'hacac;
    LUT4 mux_2169_i4_3_lut (.A(n4472), .B(n4497), .C(n19942), .Z(subOut_24__N_1369[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i4_3_lut.init = 16'hacac;
    LUT4 mux_2169_i5_3_lut (.A(n4471), .B(n4496), .C(n19942), .Z(subOut_24__N_1369[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i5_3_lut.init = 16'hacac;
    LUT4 mux_2169_i6_3_lut (.A(n4470), .B(n4495), .C(n19942), .Z(subOut_24__N_1369[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i6_3_lut.init = 16'hacac;
    LUT4 mux_2169_i7_3_lut (.A(n4469), .B(n4494), .C(n19942), .Z(subOut_24__N_1369[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i7_3_lut.init = 16'hacac;
    LUT4 mux_2169_i8_3_lut (.A(n4468), .B(n4493), .C(n19942), .Z(subOut_24__N_1369[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i8_3_lut.init = 16'hacac;
    LUT4 mux_2169_i9_3_lut (.A(n4467), .B(n4492), .C(n19942), .Z(subOut_24__N_1369[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i9_3_lut.init = 16'hacac;
    LUT4 mux_2169_i10_3_lut (.A(n4466), .B(n4491), .C(n19942), .Z(subOut_24__N_1369[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i10_3_lut.init = 16'hacac;
    LUT4 mux_2169_i11_3_lut (.A(n4465), .B(n4490), .C(n19942), .Z(subOut_24__N_1369[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i11_3_lut.init = 16'hacac;
    FD1S3AX rst_12 (.D(n21649), .CK(clkout_c), .Q(rst));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12.GSR = "DISABLED";
    GSR GSR_INST (.GSR(n22435));
    LUT4 mux_2169_i12_3_lut (.A(n4464), .B(n4489), .C(n19942), .Z(subOut_24__N_1369[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i12_3_lut.init = 16'hacac;
    LUT4 mux_2169_i13_3_lut (.A(n4463), .B(n4488), .C(n19942), .Z(subOut_24__N_1369[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i13_3_lut.init = 16'hacac;
    LUT4 mux_2169_i14_3_lut (.A(n4462), .B(n4487), .C(n19942), .Z(subOut_24__N_1369[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i14_3_lut.init = 16'hacac;
    LUT4 mux_2169_i15_3_lut (.A(n4461), .B(n4486), .C(n19942), .Z(subOut_24__N_1369[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i15_3_lut.init = 16'hacac;
    LUT4 mux_2169_i16_3_lut (.A(n4460), .B(n4485), .C(n19942), .Z(subOut_24__N_1369[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i16_3_lut.init = 16'hacac;
    LUT4 mux_2169_i17_3_lut (.A(n4459), .B(n4484), .C(n19942), .Z(subOut_24__N_1369[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i17_3_lut.init = 16'hacac;
    LUT4 mux_2169_i18_3_lut (.A(n4458), .B(n4483), .C(n19942), .Z(subOut_24__N_1369[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i18_3_lut.init = 16'hacac;
    LUT4 mux_2169_i19_3_lut (.A(n4457), .B(n4482), .C(n19942), .Z(subOut_24__N_1369[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i19_3_lut.init = 16'hacac;
    LUT4 mux_2169_i20_3_lut (.A(n4456), .B(n4481), .C(n19942), .Z(subOut_24__N_1369[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i20_3_lut.init = 16'hacac;
    LUT4 mux_2169_i21_3_lut (.A(n4455), .B(n4480), .C(n19942), .Z(subOut_24__N_1369[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i21_3_lut.init = 16'hacac;
    LUT4 mux_2169_i22_3_lut (.A(n4454), .B(n4479), .C(n19942), .Z(subOut_24__N_1369[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i22_3_lut.init = 16'hacac;
    LUT4 mux_2169_i25_3_lut (.A(n4453), .B(n4479), .C(n19942), .Z(subOut_24__N_1369[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2169_i25_3_lut.init = 16'hacac;
    LUT4 i1746_3_lut_rep_382 (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .Z(n21695)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i1746_3_lut_rep_382.init = 16'h4242;
    LUT4 i17560_2_lut_4_lut (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .D(free_m4), .Z(n3290)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i17560_2_lut_4_lut.init = 16'hffbd;
    LUT4 i1656_3_lut_rep_389 (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .Z(n21702)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i1656_3_lut_rep_389.init = 16'h4242;
    LUT4 i17562_2_lut_4_lut (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .D(free_m3), .Z(n3182)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i17562_2_lut_4_lut.init = 16'hffbd;
    COMMUTATION_U6 COM_I_M3 (.MB_m3_c_0(MB_m3_c_0), .clkout_c(clkout_c), 
            .MC_m3_c_0(MC_m3_c_0), .MA_m3_c_0(MA_m3_c_0), .LED3_c(LED3_c), 
            .enable_m3(enable_m3), .n3088(n3088), .n21705(n21705), .PWM_m3(PWM_m3), 
            .n3124(n3124), .n21703(n21703), .n19845(n19845), .n21702(n21702), 
            .free_m3(free_m3), .MA_m3_c_1(MA_m3_c_1), .n3182(n3182), .MC_m3_c_1(MC_m3_c_1), 
            .n3136(n3136), .MB_m3_c_1(MB_m3_c_1), .n3100(n3100));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(339[13:24])
    COMMUTATION_U7 COM_I_M2 (.MB_m2_c_0(MB_m2_c_0), .clkout_c(clkout_c), 
            .MC_m2_c_0(MC_m2_c_0), .MA_m2_c_0(MA_m2_c_0), .LED2_c(LED2_c), 
            .enable_m2(enable_m2), .n2980(n2980), .n21712(n21712), .PWM_m2(PWM_m2), 
            .n3016(n3016), .n21710(n21710), .n19830(n19830), .n21709(n21709), 
            .free_m2(free_m2), .MA_m2_c_1(MA_m2_c_1), .n3074(n3074), .MC_m2_c_1(MC_m2_c_1), 
            .n3028(n3028), .MB_m2_c_1(MB_m2_c_1), .n2992(n2992));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(329[13:24])
    COMMUTATION_U8 COM_I_M1 (.MB_m1_c_0(MB_m1_c_0), .clkout_c(clkout_c), 
            .MC_m1_c_0(MC_m1_c_0), .MA_m1_c_0(MA_m1_c_0), .LED1_c(LED1_c), 
            .enable_m1(enable_m1), .n2872(n2872), .n21716(n21716), .PWM_m1(PWM_m1), 
            .n2908(n2908), .n21714(n21714), .n19843(n19843), .n21713(n21713), 
            .free_m1(free_m1), .MA_m1_c_1(MA_m1_c_1), .n2966(n2966), .MC_m1_c_1(MC_m1_c_1), 
            .n2920(n2920), .MB_m1_c_1(MB_m1_c_1), .n2884(n2884));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(319[13:24])
    CLKDIV CLKDIV_I (.clkout_c(clkout_c), .clk_1mhz(clk_1mhz), .pwm_clk(pwm_clk), 
           .GND_net(GND_net), .clk_N_875(clk_N_875));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(302[14:20])
    LUT4 i1566_3_lut_rep_396 (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .Z(n21709)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i1566_3_lut_rep_396.init = 16'h4242;
    LUT4 i17564_2_lut_4_lut (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .D(free_m2), .Z(n3074)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i17564_2_lut_4_lut.init = 16'hffbd;
    LUT4 i1476_3_lut_rep_400 (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .Z(n21713)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i1476_3_lut_rep_400.init = 16'h4242;
    LUT4 i17566_2_lut_4_lut (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .D(free_m1), .Z(n2966)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i17566_2_lut_4_lut.init = 16'hffbd;
    LUT4 i2365_4_lut_rep_336 (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18836), .Z(n21649)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2365_4_lut_rep_336.init = 16'hccc8;
    LUT4 i9309_1_lut_4_lut (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18836), .Z(clkout_c_enable_362)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i9309_1_lut_4_lut.init = 16'h3337;
    HALL_U5 HALL_I_M1 (.clk_1mhz(clk_1mhz), .\speed_m1[0] (speed_m1[0]), 
            .hallsense_m1({hallsense_m1}), .clkout_c_enable_341(clkout_c_enable_341), 
            .clkout_c_enable_272(clkout_c_enable_272), .HALL_A_OUT_c_c(HALL_A_OUT_c_c), 
            .HALL_B_OUT_c_c(HALL_B_OUT_c_c), .HALL_C_OUT_c_c(HALL_C_OUT_c_c), 
            .\speed_m1[1] (speed_m1[1]), .\speed_m1[2] (speed_m1[2]), .\speed_m1[3] (speed_m1[3]), 
            .\speed_m1[4] (speed_m1[4]), .\speed_m1[5] (speed_m1[5]), .\speed_m1[6] (speed_m1[6]), 
            .\speed_m1[7] (speed_m1[7]), .\speed_m1[8] (speed_m1[8]), .\speed_m1[9] (speed_m1[9]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_m1[11] (speed_m1[11]), 
            .\speed_m1[12] (speed_m1[12]), .\speed_m1[13] (speed_m1[13]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_m1[15] (speed_m1[15]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_m1[17] (speed_m1[17]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_m1[19] (speed_m1[19]), 
            .n22430(n22430), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(316[14:18])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    AVG_SPEED AVG_SPEED_M4 (.\speed_avg_m4[0] (speed_avg_m4[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m4[0] (speed_m4[0]), .GND_net(GND_net), .\speed_avg_m4[1] (speed_avg_m4[1]), 
            .\speed_m4[1] (speed_m4[1]), .\speed_avg_m4[2] (speed_avg_m4[2]), 
            .\speed_m4[2] (speed_m4[2]), .\speed_avg_m4[3] (speed_avg_m4[3]), 
            .\speed_m4[3] (speed_m4[3]), .\speed_avg_m4[4] (speed_avg_m4[4]), 
            .\speed_m4[4] (speed_m4[4]), .\speed_avg_m4[5] (speed_avg_m4[5]), 
            .\speed_m4[5] (speed_m4[5]), .\speed_avg_m4[6] (speed_avg_m4[6]), 
            .\speed_m4[6] (speed_m4[6]), .\speed_avg_m4[7] (speed_avg_m4[7]), 
            .\speed_m4[7] (speed_m4[7]), .\speed_avg_m4[8] (speed_avg_m4[8]), 
            .\speed_m4[8] (speed_m4[8]), .\speed_avg_m4[9] (speed_avg_m4[9]), 
            .\speed_m4[9] (speed_m4[9]), .\speed_avg_m4[10] (speed_avg_m4[10]), 
            .\speed_m4[10] (speed_m4[10]), .\speed_avg_m4[11] (speed_avg_m4[11]), 
            .\speed_m4[11] (speed_m4[11]), .\speed_avg_m4[12] (speed_avg_m4[12]), 
            .\speed_m4[12] (speed_m4[12]), .\speed_avg_m4[13] (speed_avg_m4[13]), 
            .\speed_m4[13] (speed_m4[13]), .\speed_avg_m4[14] (speed_avg_m4[14]), 
            .\speed_m4[14] (speed_m4[14]), .\speed_avg_m4[15] (speed_avg_m4[15]), 
            .\speed_m4[15] (speed_m4[15]), .\speed_avg_m4[16] (speed_avg_m4[16]), 
            .\speed_m4[16] (speed_m4[16]), .\speed_avg_m4[17] (speed_avg_m4[17]), 
            .\speed_m4[17] (speed_m4[17]), .\speed_avg_m4[18] (speed_avg_m4[18]), 
            .\speed_m4[18] (speed_m4[18]), .\speed_avg_m4[19] (speed_avg_m4[19]), 
            .\speed_m4[19] (speed_m4[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(364[17:26])
    FD1P3AX start_cnt_2097__i1 (.D(n74), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i1.GSR = "DISABLED";
    SPI SPI_I (.n22435(n22435), .speed_set_m4({speed_set_m4}), .clkout_c(clkout_c), 
        .MISO_N_816(MISO_N_816), .enable_m1(enable_m1), .enable_m2(enable_m2), 
        .enable_m3(enable_m3), .enable_m4(enable_m4), .clkout_c_enable_341(clkout_c_enable_341), 
        .CS_c(CS_c), .SCK_c(SCK_c), .speed_set_m3({speed_set_m3}), .MOSI_c(MOSI_c), 
        .GND_net(GND_net), .hallsense_m1({hallsense_m1}), .dir_m1(dir_m1), 
        .n2872(n2872), .n2908(n2908), .hallsense_m2({hallsense_m2}), .dir_m2(dir_m2), 
        .n2980(n2980), .n3016(n3016), .clkout_c_enable_272(clkout_c_enable_272), 
        .hallsense_m3({hallsense_m3}), .dir_m3(dir_m3), .n3088(n3088), 
        .n3124(n3124), .rst(rst), .hallsense_m4({hallsense_m4}), .dir_m4(dir_m4), 
        .n3196(n3196), .n3232(n3232), .n5172(n5172), .speed_set_m2({speed_set_m2}), 
        .speed_set_m1({speed_set_m1}), .free_m4(free_m4), .n19826(n19826), 
        .free_m3(free_m3), .n19845(n19845), .free_m2(free_m2), .n19830(n19830), 
        .free_m1(free_m1), .n19843(n19843));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(307[10:13])
    FD1P3AX start_cnt_2097__i2 (.D(n73), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i2.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i3 (.D(n72), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i3.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i4 (.D(n71), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i4.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i5 (.D(n70), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i5.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i6 (.D(n69), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i6.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i7 (.D(n68), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i7.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i8 (.D(n67), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i8.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i9 (.D(n66), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i9.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i10 (.D(n65), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i10.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i11 (.D(n64), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i11.GSR = "DISABLED";
    FD1P3AX start_cnt_2097__i12 (.D(n63), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(start_cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i12.GSR = "DISABLED";
    FD1S3AX start_cnt_2097__i13 (.D(n10424), .CK(clkout_c), .Q(start_cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2097__i13.GSR = "DISABLED";
    AVG_SPEED_U9 AVG_SPEED_M3 (.\speed_avg_m3[0] (speed_avg_m3[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m3[0] (speed_m3[0]), .GND_net(GND_net), .\speed_avg_m3[1] (speed_avg_m3[1]), 
            .\speed_m3[1] (speed_m3[1]), .\speed_avg_m3[2] (speed_avg_m3[2]), 
            .\speed_m3[2] (speed_m3[2]), .\speed_avg_m3[3] (speed_avg_m3[3]), 
            .\speed_m3[3] (speed_m3[3]), .\speed_avg_m3[4] (speed_avg_m3[4]), 
            .\speed_m3[4] (speed_m3[4]), .\speed_avg_m3[5] (speed_avg_m3[5]), 
            .\speed_m3[5] (speed_m3[5]), .\speed_avg_m3[6] (speed_avg_m3[6]), 
            .\speed_m3[6] (speed_m3[6]), .\speed_avg_m3[7] (speed_avg_m3[7]), 
            .\speed_m3[7] (speed_m3[7]), .\speed_avg_m3[8] (speed_avg_m3[8]), 
            .\speed_m3[8] (speed_m3[8]), .\speed_avg_m3[9] (speed_avg_m3[9]), 
            .\speed_m3[9] (speed_m3[9]), .\speed_avg_m3[10] (speed_avg_m3[10]), 
            .\speed_m3[10] (speed_m3[10]), .\speed_avg_m3[11] (speed_avg_m3[11]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_avg_m3[12] (speed_avg_m3[12]), 
            .\speed_m3[12] (speed_m3[12]), .\speed_avg_m3[13] (speed_avg_m3[13]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_avg_m3[14] (speed_avg_m3[14]), 
            .\speed_m3[14] (speed_m3[14]), .\speed_avg_m3[15] (speed_avg_m3[15]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_avg_m3[16] (speed_avg_m3[16]), 
            .\speed_m3[16] (speed_m3[16]), .\speed_avg_m3[17] (speed_avg_m3[17]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_avg_m3[18] (speed_avg_m3[18]), 
            .\speed_m3[18] (speed_m3[18]), .\speed_avg_m3[19] (speed_avg_m3[19]), 
            .\speed_m3[19] (speed_m3[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(361[17:26])
    AVG_SPEED_U10 AVG_SPEED_M2 (.GND_net(GND_net), .\speed_avg_m2[0] (speed_avg_m2[0]), 
            .clk_1mhz(clk_1mhz), .\speed_m2[0] (speed_m2[0]), .\speed_avg_m2[1] (speed_avg_m2[1]), 
            .\speed_m2[1] (speed_m2[1]), .\speed_avg_m2[2] (speed_avg_m2[2]), 
            .\speed_m2[2] (speed_m2[2]), .\speed_avg_m2[3] (speed_avg_m2[3]), 
            .\speed_m2[3] (speed_m2[3]), .\speed_avg_m2[4] (speed_avg_m2[4]), 
            .\speed_m2[4] (speed_m2[4]), .\speed_avg_m2[5] (speed_avg_m2[5]), 
            .\speed_m2[5] (speed_m2[5]), .\speed_avg_m2[6] (speed_avg_m2[6]), 
            .\speed_m2[6] (speed_m2[6]), .\speed_avg_m2[7] (speed_avg_m2[7]), 
            .\speed_m2[7] (speed_m2[7]), .\speed_avg_m2[8] (speed_avg_m2[8]), 
            .\speed_m2[8] (speed_m2[8]), .\speed_avg_m2[9] (speed_avg_m2[9]), 
            .\speed_m2[9] (speed_m2[9]), .\speed_avg_m2[10] (speed_avg_m2[10]), 
            .\speed_m2[10] (speed_m2[10]), .\speed_avg_m2[11] (speed_avg_m2[11]), 
            .\speed_m2[11] (speed_m2[11]), .\speed_avg_m2[12] (speed_avg_m2[12]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_avg_m2[13] (speed_avg_m2[13]), 
            .\speed_m2[13] (speed_m2[13]), .\speed_avg_m2[14] (speed_avg_m2[14]), 
            .\speed_m2[14] (speed_m2[14]), .\speed_avg_m2[15] (speed_avg_m2[15]), 
            .\speed_m2[15] (speed_m2[15]), .\speed_avg_m2[16] (speed_avg_m2[16]), 
            .\speed_m2[16] (speed_m2[16]), .\speed_avg_m2[17] (speed_avg_m2[17]), 
            .\speed_m2[17] (speed_m2[17]), .\speed_avg_m2[18] (speed_avg_m2[18]), 
            .\speed_m2[18] (speed_m2[18]), .\speed_avg_m2[19] (speed_avg_m2[19]), 
            .\speed_m2[19] (speed_m2[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(358[17:26])
    AVG_SPEED_U11 AVG_SPEED_M1 (.GND_net(GND_net), .\speed_avg_m1[0] (speed_avg_m1[0]), 
            .clk_1mhz(clk_1mhz), .\speed_m1[0] (speed_m1[0]), .\speed_avg_m1[1] (speed_avg_m1[1]), 
            .\speed_m1[1] (speed_m1[1]), .\speed_avg_m1[2] (speed_avg_m1[2]), 
            .\speed_m1[2] (speed_m1[2]), .\speed_avg_m1[3] (speed_avg_m1[3]), 
            .\speed_m1[3] (speed_m1[3]), .\speed_avg_m1[4] (speed_avg_m1[4]), 
            .\speed_m1[4] (speed_m1[4]), .\speed_avg_m1[5] (speed_avg_m1[5]), 
            .\speed_m1[5] (speed_m1[5]), .\speed_avg_m1[6] (speed_avg_m1[6]), 
            .\speed_m1[6] (speed_m1[6]), .\speed_avg_m1[7] (speed_avg_m1[7]), 
            .\speed_m1[7] (speed_m1[7]), .\speed_avg_m1[8] (speed_avg_m1[8]), 
            .\speed_m1[8] (speed_m1[8]), .\speed_avg_m1[9] (speed_avg_m1[9]), 
            .\speed_m1[9] (speed_m1[9]), .\speed_avg_m1[10] (speed_avg_m1[10]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_avg_m1[11] (speed_avg_m1[11]), 
            .\speed_m1[11] (speed_m1[11]), .\speed_avg_m1[12] (speed_avg_m1[12]), 
            .\speed_m1[12] (speed_m1[12]), .\speed_avg_m1[13] (speed_avg_m1[13]), 
            .\speed_m1[13] (speed_m1[13]), .\speed_avg_m1[14] (speed_avg_m1[14]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_avg_m1[15] (speed_avg_m1[15]), 
            .\speed_m1[15] (speed_m1[15]), .\speed_avg_m1[16] (speed_avg_m1[16]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_avg_m1[17] (speed_avg_m1[17]), 
            .\speed_m1[17] (speed_m1[17]), .\speed_avg_m1[18] (speed_avg_m1[18]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_avg_m1[19] (speed_avg_m1[19]), 
            .\speed_m1[19] (speed_m1[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(355[17:26])
    HALL_U3 HALL_I_M3 (.clk_1mhz(clk_1mhz), .n22430(n22430), .\speed_m3[0] (speed_m3[0]), 
            .hallsense_m3({hallsense_m3}), .clkout_c_enable_341(clkout_c_enable_341), 
            .H_A_m3_c(H_A_m3_c), .H_B_m3_c(H_B_m3_c), .H_C_m3_c(H_C_m3_c), 
            .\speed_m3[1] (speed_m3[1]), .\speed_m3[2] (speed_m3[2]), .\speed_m3[3] (speed_m3[3]), 
            .\speed_m3[4] (speed_m3[4]), .\speed_m3[5] (speed_m3[5]), .\speed_m3[6] (speed_m3[6]), 
            .\speed_m3[7] (speed_m3[7]), .\speed_m3[8] (speed_m3[8]), .\speed_m3[9] (speed_m3[9]), 
            .\speed_m3[10] (speed_m3[10]), .\speed_m3[11] (speed_m3[11]), 
            .\speed_m3[12] (speed_m3[12]), .\speed_m3[13] (speed_m3[13]), 
            .\speed_m3[14] (speed_m3[14]), .\speed_m3[15] (speed_m3[15]), 
            .\speed_m3[16] (speed_m3[16]), .\speed_m3[17] (speed_m3[17]), 
            .\speed_m3[18] (speed_m3[18]), .\speed_m3[19] (speed_m3[19]), 
            .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(336[14:18])
    FD1S3AX rst_12_rep_428 (.D(n21649), .CK(clkout_c), .Q(clkout_c_enable_341));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12_rep_428.GSR = "DISABLED";
    PWMGENERATOR_U1 PWM_I_M2 (.PWM_m2(PWM_m2), .pwm_clk(pwm_clk), .free_m2(free_m2), 
            .clkout_c_enable_341(clkout_c_enable_341), .PWMdut_m2({PWMdut_m2}), 
            .GND_net(GND_net), .hallsense_m2({hallsense_m2}), .n21710(n21710), 
            .enable_m2(enable_m2), .n3028(n3028), .n21712(n21712), .n2992(n2992));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(332[13:25])
    COMMUTATION COM_I_M4 (.MB_m4_c_0(MB_m4_c_0), .clkout_c(clkout_c), .MC_m4_c_0(MC_m4_c_0), 
            .MA_m4_c_0(MA_m4_c_0), .LED4_c(LED4_c), .enable_m4(enable_m4), 
            .n3196(n3196), .n21700(n21700), .PWM_m4(PWM_m4), .n3232(n3232), 
            .n21696(n21696), .n19826(n19826), .n21695(n21695), .free_m4(free_m4), 
            .MA_m4_c_1(MA_m4_c_1), .n3290(n3290), .MC_m4_c_1(MC_m4_c_1), 
            .n3244(n3244), .MB_m4_c_1(MB_m4_c_1), .n3208(n3208));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(349[13:24])
    PWMGENERATOR_U2 PWM_I_M1 (.PWM_m1(PWM_m1), .pwm_clk(pwm_clk), .free_m1(free_m1), 
            .clkout_c_enable_341(clkout_c_enable_341), .PWMdut_m1({PWMdut_m1}), 
            .GND_net(GND_net), .hallsense_m1({hallsense_m1}), .n21714(n21714), 
            .enable_m1(enable_m1), .n2920(n2920), .n21716(n21716), .n2884(n2884));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(322[13:25])
    PWMGENERATOR_U0 PWM_I_M3 (.PWM_m3(PWM_m3), .pwm_clk(pwm_clk), .free_m3(free_m3), 
            .clkout_c_enable_341(clkout_c_enable_341), .PWMdut_m3({PWMdut_m3}), 
            .GND_net(GND_net), .hallsense_m3({hallsense_m3}), .n21703(n21703), 
            .enable_m3(enable_m3), .n3136(n3136), .n21705(n21705), .n3100(n3100));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(342[13:25])
    HALL_U4 HALL_I_M2 (.clk_1mhz(clk_1mhz), .\speed_m2[0] (speed_m2[0]), 
            .hallsense_m2({hallsense_m2}), .rst(rst), .H_B_m2_c(H_B_m2_c), 
            .clkout_c_enable_272(clkout_c_enable_272), .H_A_m2_c(H_A_m2_c), 
            .clkout_c_enable_341(clkout_c_enable_341), .H_C_m2_c(H_C_m2_c), 
            .\speed_m2[1] (speed_m2[1]), .\speed_m2[2] (speed_m2[2]), .\speed_m2[3] (speed_m2[3]), 
            .\speed_m2[4] (speed_m2[4]), .\speed_m2[5] (speed_m2[5]), .\speed_m2[6] (speed_m2[6]), 
            .\speed_m2[7] (speed_m2[7]), .\speed_m2[8] (speed_m2[8]), .\speed_m2[9] (speed_m2[9]), 
            .\speed_m2[10] (speed_m2[10]), .\speed_m2[11] (speed_m2[11]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_m2[13] (speed_m2[13]), 
            .\speed_m2[14] (speed_m2[14]), .\speed_m2[15] (speed_m2[15]), 
            .\speed_m2[16] (speed_m2[16]), .\speed_m2[17] (speed_m2[17]), 
            .\speed_m2[18] (speed_m2[18]), .\speed_m2[19] (speed_m2[19]), 
            .GND_net(GND_net), .n22430(n22430));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(326[14:18])
    \PID(16000000,160000000,10000000)  PID_I (.GND_net(GND_net), .n4466(n4466), 
            .n4465(n4465), .speed_set_m3({speed_set_m3}), .speed_set_m4({speed_set_m4}), 
            .clk_N_875(clk_N_875), .n4468(n4468), .n4467(n4467), .n4470(n4470), 
            .n4469(n4469), .\subOut_24__N_1369[0] (subOut_24__N_1369[0]), 
            .speed_set_m2({speed_set_m2}), .PWMdut_m2({PWMdut_m2}), .speed_set_m1({speed_set_m1}), 
            .\speed_avg_m3[12] (speed_avg_m3[12]), .\speed_avg_m2[12] (speed_avg_m2[12]), 
            .\speed_avg_m3[9] (speed_avg_m3[9]), .\speed_avg_m2[9] (speed_avg_m2[9]), 
            .\speed_avg_m3[8] (speed_avg_m3[8]), .\speed_avg_m2[8] (speed_avg_m2[8]), 
            .\speed_avg_m3[7] (speed_avg_m3[7]), .\speed_avg_m2[7] (speed_avg_m2[7]), 
            .\speed_avg_m3[3] (speed_avg_m3[3]), .\speed_avg_m2[3] (speed_avg_m2[3]), 
            .\speed_avg_m4[19] (speed_avg_m4[19]), .\speed_avg_m3[19] (speed_avg_m3[19]), 
            .\speed_avg_m4[18] (speed_avg_m4[18]), .\speed_avg_m3[18] (speed_avg_m3[18]), 
            .\speed_avg_m4[17] (speed_avg_m4[17]), .\speed_avg_m3[17] (speed_avg_m3[17]), 
            .\speed_avg_m4[16] (speed_avg_m4[16]), .\speed_avg_m3[16] (speed_avg_m3[16]), 
            .\speed_avg_m4[15] (speed_avg_m4[15]), .\speed_avg_m3[15] (speed_avg_m3[15]), 
            .\speed_avg_m4[14] (speed_avg_m4[14]), .\speed_avg_m3[14] (speed_avg_m3[14]), 
            .\speed_avg_m4[13] (speed_avg_m4[13]), .\speed_avg_m3[13] (speed_avg_m3[13]), 
            .\speed_avg_m4[11] (speed_avg_m4[11]), .\speed_avg_m3[11] (speed_avg_m3[11]), 
            .\speed_avg_m4[10] (speed_avg_m4[10]), .\speed_avg_m3[10] (speed_avg_m3[10]), 
            .\speed_avg_m4[6] (speed_avg_m4[6]), .\speed_avg_m3[6] (speed_avg_m3[6]), 
            .dir_m2(dir_m2), .dir_m3(dir_m3), .dir_m1(dir_m1), .dir_m4(dir_m4), 
            .\speed_avg_m4[5] (speed_avg_m4[5]), .\speed_avg_m3[5] (speed_avg_m3[5]), 
            .\speed_avg_m4[4] (speed_avg_m4[4]), .\speed_avg_m3[4] (speed_avg_m3[4]), 
            .n4472(n4472), .n4471(n4471), .\speed_avg_m4[2] (speed_avg_m4[2]), 
            .\speed_avg_m3[2] (speed_avg_m3[2]), .\speed_avg_m4[1] (speed_avg_m4[1]), 
            .\speed_avg_m3[1] (speed_avg_m3[1]), .\speed_avg_m4[0] (speed_avg_m4[0]), 
            .\speed_avg_m3[0] (speed_avg_m3[0]), .VCC_net(VCC_net), .\speed_avg_m1[12] (speed_avg_m1[12]), 
            .\speed_avg_m1[9] (speed_avg_m1[9]), .\speed_avg_m1[8] (speed_avg_m1[8]), 
            .n4474(n4474), .n4473(n4473), .\speed_avg_m1[7] (speed_avg_m1[7]), 
            .\speed_avg_m1[3] (speed_avg_m1[3]), .\speed_avg_m1[19] (speed_avg_m1[19]), 
            .\speed_avg_m2[19] (speed_avg_m2[19]), .\speed_avg_m1[18] (speed_avg_m1[18]), 
            .\speed_avg_m2[18] (speed_avg_m2[18]), .\speed_avg_m1[17] (speed_avg_m1[17]), 
            .\speed_avg_m2[17] (speed_avg_m2[17]), .\speed_avg_m1[16] (speed_avg_m1[16]), 
            .\speed_avg_m2[16] (speed_avg_m2[16]), .\speed_avg_m1[15] (speed_avg_m1[15]), 
            .\speed_avg_m2[15] (speed_avg_m2[15]), .\speed_avg_m1[14] (speed_avg_m1[14]), 
            .\speed_avg_m2[14] (speed_avg_m2[14]), .\speed_avg_m1[13] (speed_avg_m1[13]), 
            .\speed_avg_m2[13] (speed_avg_m2[13]), .\speed_avg_m1[11] (speed_avg_m1[11]), 
            .\speed_avg_m2[11] (speed_avg_m2[11]), .\speed_avg_m1[10] (speed_avg_m1[10]), 
            .\speed_avg_m2[10] (speed_avg_m2[10]), .\speed_avg_m1[6] (speed_avg_m1[6]), 
            .\speed_avg_m2[6] (speed_avg_m2[6]), .\speed_avg_m1[5] (speed_avg_m1[5]), 
            .\speed_avg_m2[5] (speed_avg_m2[5]), .\speed_avg_m1[4] (speed_avg_m1[4]), 
            .\speed_avg_m2[4] (speed_avg_m2[4]), .\speed_avg_m1[2] (speed_avg_m1[2]), 
            .\speed_avg_m2[2] (speed_avg_m2[2]), .\speed_avg_m1[1] (speed_avg_m1[1]), 
            .\speed_avg_m2[1] (speed_avg_m2[1]), .\speed_avg_m1[0] (speed_avg_m1[0]), 
            .\speed_avg_m2[0] (speed_avg_m2[0]), .n4475(n4475), .\subOut_24__N_1369[1] (subOut_24__N_1369[1]), 
            .\subOut_24__N_1369[2] (subOut_24__N_1369[2]), .\subOut_24__N_1369[3] (subOut_24__N_1369[3]), 
            .\subOut_24__N_1369[4] (subOut_24__N_1369[4]), .\subOut_24__N_1369[5] (subOut_24__N_1369[5]), 
            .\subOut_24__N_1369[6] (subOut_24__N_1369[6]), .\subOut_24__N_1369[7] (subOut_24__N_1369[7]), 
            .\subOut_24__N_1369[8] (subOut_24__N_1369[8]), .\subOut_24__N_1369[9] (subOut_24__N_1369[9]), 
            .\subOut_24__N_1369[10] (subOut_24__N_1369[10]), .\subOut_24__N_1369[11] (subOut_24__N_1369[11]), 
            .\subOut_24__N_1369[12] (subOut_24__N_1369[12]), .\subOut_24__N_1369[13] (subOut_24__N_1369[13]), 
            .\subOut_24__N_1369[14] (subOut_24__N_1369[14]), .\subOut_24__N_1369[15] (subOut_24__N_1369[15]), 
            .\subOut_24__N_1369[16] (subOut_24__N_1369[16]), .\subOut_24__N_1369[17] (subOut_24__N_1369[17]), 
            .\subOut_24__N_1369[18] (subOut_24__N_1369[18]), .\subOut_24__N_1369[19] (subOut_24__N_1369[19]), 
            .\subOut_24__N_1369[20] (subOut_24__N_1369[20]), .\subOut_24__N_1369[21] (subOut_24__N_1369[21]), 
            .\subOut_24__N_1369[24] (subOut_24__N_1369[24]), .n19942(n19942), 
            .n22435(n22435), .PWMdut_m1({PWMdut_m1}), .\speed_avg_m4[12] (speed_avg_m4[12]), 
            .\speed_avg_m4[9] (speed_avg_m4[9]), .\speed_avg_m4[8] (speed_avg_m4[8]), 
            .\speed_avg_m4[7] (speed_avg_m4[7]), .\speed_avg_m4[3] (speed_avg_m4[3]), 
            .n4479(n4479), .n4481(n4481), .n4480(n4480), .n4483(n4483), 
            .n4482(n4482), .PWMdut_m4({PWMdut_m4}), .n4485(n4485), .n4484(n4484), 
            .PWMdut_m3({PWMdut_m3}), .n4487(n4487), .n4486(n4486), .n4489(n4489), 
            .n4488(n4488), .n4491(n4491), .n4490(n4490), .n4493(n4493), 
            .n4492(n4492), .n4495(n4495), .n4494(n4494), .n4497(n4497), 
            .n4496(n4496), .n4499(n4499), .n4498(n4498), .n4500(n4500), 
            .n4454(n4454), .n4453(n4453), .n4456(n4456), .n4455(n4455), 
            .n4458(n4458), .n4457(n4457), .n4460(n4460), .n4459(n4459), 
            .n4462(n4462), .n4461(n4461), .n4464(n4464), .n4463(n4463));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(311[10:13])
    FD1S3AX rst_12_rep_427 (.D(n21649), .CK(clkout_c), .Q(clkout_c_enable_272));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12_rep_427.GSR = "DISABLED";
    PWMGENERATOR PWM_I_M4 (.pwm_clk(pwm_clk), .PWM_m4(PWM_m4), .free_m4(free_m4), 
            .clkout_c_enable_341(clkout_c_enable_341), .PWMdut_m4({PWMdut_m4}), 
            .GND_net(GND_net), .hallsense_m4({hallsense_m4}), .n21696(n21696), 
            .enable_m4(enable_m4), .n3244(n3244), .n21700(n21700), .n3208(n3208));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(352[13:25])
    HALL HALL_I_M4 (.clk_1mhz(clk_1mhz), .\speed_m4[0] (speed_m4[0]), .hallsense_m4({hallsense_m4}), 
         .clkout_c_enable_272(clkout_c_enable_272), .clkout_c_enable_341(clkout_c_enable_341), 
         .H_A_m4_c(H_A_m4_c), .H_B_m4_c(H_B_m4_c), .H_C_m4_c(H_C_m4_c), 
         .\speed_m4[1] (speed_m4[1]), .\speed_m4[2] (speed_m4[2]), .\speed_m4[3] (speed_m4[3]), 
         .\speed_m4[4] (speed_m4[4]), .\speed_m4[5] (speed_m4[5]), .\speed_m4[6] (speed_m4[6]), 
         .\speed_m4[7] (speed_m4[7]), .\speed_m4[8] (speed_m4[8]), .\speed_m4[9] (speed_m4[9]), 
         .\speed_m4[10] (speed_m4[10]), .\speed_m4[11] (speed_m4[11]), .\speed_m4[12] (speed_m4[12]), 
         .\speed_m4[13] (speed_m4[13]), .\speed_m4[14] (speed_m4[14]), .\speed_m4[15] (speed_m4[15]), 
         .\speed_m4[16] (speed_m4[16]), .\speed_m4[17] (speed_m4[17]), .\speed_m4[18] (speed_m4[18]), 
         .\speed_m4[19] (speed_m4[19]), .GND_net(GND_net), .n22430(n22430));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(346[14:18])
    
endmodule
//
// Verilog Description of module COMMUTATION_U6
//

module COMMUTATION_U6 (MB_m3_c_0, clkout_c, MC_m3_c_0, MA_m3_c_0, LED3_c, 
            enable_m3, n3088, n21705, PWM_m3, n3124, n21703, n19845, 
            n21702, free_m3, MA_m3_c_1, n3182, MC_m3_c_1, n3136, 
            MB_m3_c_1, n3100);
    output MB_m3_c_0;
    input clkout_c;
    output MC_m3_c_0;
    output MA_m3_c_0;
    output LED3_c;
    input enable_m3;
    input n3088;
    input n21705;
    input PWM_m3;
    input n3124;
    input n21703;
    input n19845;
    input n21702;
    input free_m3;
    output MA_m3_c_1;
    input n3182;
    output MC_m3_c_1;
    input n3136;
    output MB_m3_c_1;
    input n3100;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_2151, n18970, n18969, n19846, n14107;
    
    FD1S3IX MospairB_i1 (.D(n18970), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MB_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18969), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MC_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19846), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MA_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14107), .CK(clkout_c), .PD(led1_N_2151), .Q(LED3_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10634_1_lut (.A(enable_m3), .Z(led1_N_2151)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10634_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3088), .B(n21705), .C(PWM_m3), .Z(n18970)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_201 (.A(n3124), .B(n21703), .C(PWM_m3), .Z(n18969)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_201.init = 16'hbfbf;
    LUT4 i17576_3_lut (.A(n19845), .B(PWM_m3), .C(n21702), .Z(n19846)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17576_3_lut.init = 16'hbfbf;
    LUT4 i11520_2_lut (.A(free_m3), .B(LED3_c), .Z(n14107)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11520_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n3182), .CK(clkout_c), .CD(n19845), .Q(MA_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3124), .CK(clkout_c), .CD(n3136), .Q(MC_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3088), .CK(clkout_c), .CD(n3100), .Q(MB_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION_U7
//

module COMMUTATION_U7 (MB_m2_c_0, clkout_c, MC_m2_c_0, MA_m2_c_0, LED2_c, 
            enable_m2, n2980, n21712, PWM_m2, n3016, n21710, n19830, 
            n21709, free_m2, MA_m2_c_1, n3074, MC_m2_c_1, n3028, 
            MB_m2_c_1, n2992);
    output MB_m2_c_0;
    input clkout_c;
    output MC_m2_c_0;
    output MA_m2_c_0;
    output LED2_c;
    input enable_m2;
    input n2980;
    input n21712;
    input PWM_m2;
    input n3016;
    input n21710;
    input n19830;
    input n21709;
    input free_m2;
    output MA_m2_c_1;
    input n3074;
    output MC_m2_c_1;
    input n3028;
    output MB_m2_c_1;
    input n2992;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_2151, n18972, n18971, n19831, n14109;
    
    FD1S3IX MospairB_i1 (.D(n18972), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MB_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18971), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MC_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19831), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MA_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14109), .CK(clkout_c), .PD(led1_N_2151), .Q(LED2_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10633_1_lut (.A(enable_m2), .Z(led1_N_2151)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10633_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2980), .B(n21712), .C(PWM_m2), .Z(n18972)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_200 (.A(n3016), .B(n21710), .C(PWM_m2), .Z(n18971)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_200.init = 16'hbfbf;
    LUT4 i17578_3_lut (.A(n19830), .B(PWM_m2), .C(n21709), .Z(n19831)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17578_3_lut.init = 16'hbfbf;
    LUT4 i11522_2_lut (.A(free_m2), .B(LED2_c), .Z(n14109)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11522_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n3074), .CK(clkout_c), .CD(n19830), .Q(MA_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3016), .CK(clkout_c), .CD(n3028), .Q(MC_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2980), .CK(clkout_c), .CD(n2992), .Q(MB_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION_U8
//

module COMMUTATION_U8 (MB_m1_c_0, clkout_c, MC_m1_c_0, MA_m1_c_0, LED1_c, 
            enable_m1, n2872, n21716, PWM_m1, n2908, n21714, n19843, 
            n21713, free_m1, MA_m1_c_1, n2966, MC_m1_c_1, n2920, 
            MB_m1_c_1, n2884);
    output MB_m1_c_0;
    input clkout_c;
    output MC_m1_c_0;
    output MA_m1_c_0;
    output LED1_c;
    input enable_m1;
    input n2872;
    input n21716;
    input PWM_m1;
    input n2908;
    input n21714;
    input n19843;
    input n21713;
    input free_m1;
    output MA_m1_c_1;
    input n2966;
    output MC_m1_c_1;
    input n2920;
    output MB_m1_c_1;
    input n2884;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_2151, n18974, n18973, n19844, n14111;
    
    FD1S3IX MospairB_i1 (.D(n18974), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MB_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18973), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MC_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19844), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MA_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14111), .CK(clkout_c), .PD(led1_N_2151), .Q(LED1_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10630_1_lut (.A(enable_m1), .Z(led1_N_2151)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10630_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2872), .B(n21716), .C(PWM_m1), .Z(n18974)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_199 (.A(n2908), .B(n21714), .C(PWM_m1), .Z(n18973)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_199.init = 16'hbfbf;
    LUT4 i17585_3_lut (.A(n19843), .B(PWM_m1), .C(n21713), .Z(n19844)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17585_3_lut.init = 16'hbfbf;
    LUT4 i11524_2_lut (.A(free_m1), .B(LED1_c), .Z(n14111)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11524_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n2966), .CK(clkout_c), .CD(n19843), .Q(MA_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n2908), .CK(clkout_c), .CD(n2920), .Q(MC_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2872), .CK(clkout_c), .CD(n2884), .Q(MB_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module CLKDIV
//

module CLKDIV (clkout_c, clk_1mhz, pwm_clk, GND_net, clk_N_875);
    input clkout_c;
    output clk_1mhz;
    output pwm_clk;
    input GND_net;
    output clk_N_875;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    wire pi_clk /* synthesis is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(89[9:15])
    wire clk_N_875 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    
    wire mhz_buf, mhz_buf_N_68, pi_buf, pi_buf_N_69, pwm_buf, pwm_buf_N_67, 
        n14145, n20148;
    wire [11:0]cntpi;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(42[8:13])
    
    wire n20142, n14146;
    wire [4:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(41[8:13])
    wire [4:0]n25;
    
    wire n21701, n20104;
    wire [8:0]n41;
    
    wire n18531, n18530, n18529, n18528;
    
    FD1S3AX mhz_buf_29 (.D(mhz_buf_N_68), .CK(clkout_c), .Q(mhz_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam mhz_buf_29.GSR = "DISABLED";
    FD1S3AX pi_buf_30 (.D(pi_buf_N_69), .CK(clkout_c), .Q(pi_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pi_buf_30.GSR = "DISABLED";
    FD1S3AX pwm_buf_32 (.D(pwm_buf_N_67), .CK(clkout_c), .Q(pwm_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pwm_buf_32.GSR = "DISABLED";
    FD1S3AX clk_1mhz_33 (.D(mhz_buf), .CK(clkout_c), .Q(clk_1mhz)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam clk_1mhz_33.GSR = "DISABLED";
    FD1S3AX pwm_clk_34 (.D(pwm_buf), .CK(clkout_c), .Q(pwm_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pwm_clk_34.GSR = "DISABLED";
    FD1S3AX pi_clk_35 (.D(pi_buf), .CK(clkout_c), .Q(pi_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pi_clk_35.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(pi_buf), .B(n14145), .Z(pi_buf_N_69)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    LUT4 i17478_4_lut (.A(n20148), .B(cntpi[2]), .C(n20142), .D(cntpi[7]), 
         .Z(n14145)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(66[5:16])
    defparam i17478_4_lut.init = 16'h0020;
    LUT4 i16750_3_lut (.A(cntpi[3]), .B(cntpi[8]), .C(cntpi[1]), .Z(n20148)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16750_3_lut.init = 16'h8080;
    LUT4 i16744_4_lut (.A(cntpi[0]), .B(cntpi[6]), .C(cntpi[5]), .D(cntpi[4]), 
         .Z(n20142)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16744_4_lut.init = 16'h8000;
    LUT4 pwm_buf_I_0_1_lut (.A(pwm_buf), .Z(pwm_buf_N_67)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(73[14:25])
    defparam pwm_buf_I_0_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_198 (.A(mhz_buf), .B(n14146), .Z(mhz_buf_N_68)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_198.init = 16'h6666;
    LUT4 i15399_2_lut (.A(count[1]), .B(count[0]), .Z(n25[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15399_2_lut.init = 16'h6666;
    LUT4 i15420_3_lut_4_lut (.A(count[2]), .B(n21701), .C(count[3]), .D(count[4]), 
         .Z(n25[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15420_3_lut_4_lut.init = 16'h7f80;
    LUT4 i17482_4_lut (.A(count[3]), .B(count[2]), .C(count[0]), .D(n20104), 
         .Z(n14146)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(61[5:15])
    defparam i17482_4_lut.init = 16'h1000;
    LUT4 i16706_2_lut (.A(count[1]), .B(count[4]), .Z(n20104)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16706_2_lut.init = 16'h8888;
    LUT4 i15397_1_lut (.A(count[0]), .Z(n25[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15397_1_lut.init = 16'h5555;
    FD1S3IX cntpi_2099_2100__i2 (.D(n41[1]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i2.GSR = "DISABLED";
    CCU2D cntpi_2099_2100_add_4_9 (.A0(cntpi[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18531), .S0(n41[7]), .S1(n41[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100_add_4_9.INIT0 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_9.INIT1 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_9.INJECT1_0 = "NO";
    defparam cntpi_2099_2100_add_4_9.INJECT1_1 = "NO";
    CCU2D cntpi_2099_2100_add_4_7 (.A0(cntpi[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18530), .COUT(n18531), .S0(n41[5]), .S1(n41[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100_add_4_7.INIT0 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_7.INIT1 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_7.INJECT1_0 = "NO";
    defparam cntpi_2099_2100_add_4_7.INJECT1_1 = "NO";
    CCU2D cntpi_2099_2100_add_4_5 (.A0(cntpi[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18529), .COUT(n18530), .S0(n41[3]), .S1(n41[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100_add_4_5.INIT0 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_5.INIT1 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_5.INJECT1_0 = "NO";
    defparam cntpi_2099_2100_add_4_5.INJECT1_1 = "NO";
    CCU2D cntpi_2099_2100_add_4_3 (.A0(cntpi[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18528), .COUT(n18529), .S0(n41[1]), .S1(n41[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100_add_4_3.INIT0 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_3.INIT1 = 16'hfaaa;
    defparam cntpi_2099_2100_add_4_3.INJECT1_0 = "NO";
    defparam cntpi_2099_2100_add_4_3.INJECT1_1 = "NO";
    CCU2D cntpi_2099_2100_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18528), .S1(n41[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100_add_4_1.INIT0 = 16'hF000;
    defparam cntpi_2099_2100_add_4_1.INIT1 = 16'h0555;
    defparam cntpi_2099_2100_add_4_1.INJECT1_0 = "NO";
    defparam cntpi_2099_2100_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2098__i0 (.D(n25[0]), .CK(clkout_c), .CD(n14146), .Q(count[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2098__i0.GSR = "DISABLED";
    LUT4 i15402_2_lut_rep_388 (.A(count[1]), .B(count[0]), .Z(n21701)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15402_2_lut_rep_388.init = 16'h8888;
    LUT4 i15406_2_lut_3_lut (.A(count[1]), .B(count[0]), .C(count[2]), 
         .Z(n25[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15406_2_lut_3_lut.init = 16'h7878;
    LUT4 i15413_2_lut_3_lut_4_lut (.A(count[1]), .B(count[0]), .C(count[3]), 
         .D(count[2]), .Z(n25[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15413_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1S3IX cntpi_2099_2100__i1 (.D(n41[0]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i1.GSR = "DISABLED";
    INV i17831 (.A(pi_clk), .Z(clk_N_875));
    FD1S3IX cntpi_2099_2100__i3 (.D(n41[2]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i3.GSR = "DISABLED";
    FD1S3IX cntpi_2099_2100__i4 (.D(n41[3]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i4.GSR = "DISABLED";
    FD1S3IX cntpi_2099_2100__i5 (.D(n41[4]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i5.GSR = "DISABLED";
    FD1S3IX cntpi_2099_2100__i6 (.D(n41[5]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i6.GSR = "DISABLED";
    FD1S3IX cntpi_2099_2100__i7 (.D(n41[6]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i7.GSR = "DISABLED";
    FD1S3IX cntpi_2099_2100__i8 (.D(n41[7]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i8.GSR = "DISABLED";
    FD1S3IX cntpi_2099_2100__i9 (.D(n41[8]), .CK(clkout_c), .CD(n14145), 
            .Q(cntpi[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2099_2100__i9.GSR = "DISABLED";
    FD1S3IX count_2098__i1 (.D(n25[1]), .CK(clkout_c), .CD(n14146), .Q(count[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2098__i1.GSR = "DISABLED";
    FD1S3IX count_2098__i2 (.D(n25[2]), .CK(clkout_c), .CD(n14146), .Q(count[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2098__i2.GSR = "DISABLED";
    FD1S3IX count_2098__i3 (.D(n25[3]), .CK(clkout_c), .CD(n14146), .Q(count[3]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2098__i3.GSR = "DISABLED";
    FD1S3IX count_2098__i4 (.D(n25[4]), .CK(clkout_c), .CD(n14146), .Q(count[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2098__i4.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module HALL_U5
//

module HALL_U5 (clk_1mhz, \speed_m1[0] , hallsense_m1, clkout_c_enable_341, 
            clkout_c_enable_272, HALL_A_OUT_c_c, HALL_B_OUT_c_c, HALL_C_OUT_c_c, 
            \speed_m1[1] , \speed_m1[2] , \speed_m1[3] , \speed_m1[4] , 
            \speed_m1[5] , \speed_m1[6] , \speed_m1[7] , \speed_m1[8] , 
            \speed_m1[9] , \speed_m1[10] , \speed_m1[11] , \speed_m1[12] , 
            \speed_m1[13] , \speed_m1[14] , \speed_m1[15] , \speed_m1[16] , 
            \speed_m1[17] , \speed_m1[18] , \speed_m1[19] , n22430, 
            GND_net);
    input clk_1mhz;
    output \speed_m1[0] ;
    output [2:0]hallsense_m1;
    input clkout_c_enable_341;
    input clkout_c_enable_272;
    input HALL_A_OUT_c_c;
    input HALL_B_OUT_c_c;
    input HALL_C_OUT_c_c;
    output \speed_m1[1] ;
    output \speed_m1[2] ;
    output \speed_m1[3] ;
    output \speed_m1[4] ;
    output \speed_m1[5] ;
    output \speed_m1[6] ;
    output \speed_m1[7] ;
    output \speed_m1[8] ;
    output \speed_m1[9] ;
    output \speed_m1[10] ;
    output \speed_m1[11] ;
    output \speed_m1[12] ;
    output \speed_m1[13] ;
    output \speed_m1[14] ;
    output \speed_m1[15] ;
    output \speed_m1[16] ;
    output \speed_m1[17] ;
    output \speed_m1[18] ;
    output \speed_m1[19] ;
    input n22430;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_70;
    wire [19:0]count_19__N_2067;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21661, n11471, n11469, stable_counting, stable_counting_N_2129, 
        n19815, n20042, n20184, n20160;
    wire [19:0]speedt_19__N_2047;
    
    wire hall3_lat;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n20156, n20048, n4585, n19937, n21654, n19814, n21683, 
        n21644, n4, n21640;
    wire [6:0]n63;
    
    wire hall1_old, hall1_lat, hall2_old, hall2_lat, hall3_old, n4_adj_2426, 
        n12, n19075, n20034, clk_1mhz_enable_187, n19, n24, n20, 
        n22, n16, n21682, n21724, n21651, n14402, n18462, n18461, 
        n18460, n18459, n18458, n18457, n18456, n18455, n18454, 
        n18453;
    
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2067[0]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    LUT4 i2403_2_lut_rep_348_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21661)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2403_2_lut_rep_348_3_lut_4_lut.init = 16'h8000;
    LUT4 i11515_4_lut (.A(n11471), .B(n11469), .C(stable_counting), .D(stable_counting_N_2129), 
         .Z(clk_1mhz_enable_70)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11515_4_lut.init = 16'hcaea;
    LUT4 i1_4_lut (.A(n19815), .B(n20042), .C(n20184), .D(n20160), .Z(n11471)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0002;
    FD1P3AX speed__i1 (.D(speedt_19__N_2047[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    LUT4 i16645_2_lut (.A(count[18]), .B(count[1]), .Z(n20042)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16645_2_lut.init = 16'heeee;
    LUT4 i16786_4_lut (.A(count[7]), .B(n20156), .C(n20048), .D(count[15]), 
         .Z(n20184)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16786_4_lut.init = 16'hfffe;
    LUT4 i16762_3_lut (.A(count[5]), .B(count[17]), .C(count[16]), .Z(n20160)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16762_3_lut.init = 16'hfefe;
    LUT4 i16758_4_lut (.A(count[11]), .B(count[12]), .C(count[4]), .D(count[6]), 
         .Z(n20156)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16758_4_lut.init = 16'hfffe;
    FD1S3IX count__i0 (.D(count_19__N_2067[0]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    LUT4 i16651_2_lut (.A(count[19]), .B(count[14]), .Z(n20048)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16651_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(n19937), .B(stable_count[0]), .C(n21654), .D(n19814), 
         .Z(n11469)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    LUT4 i2415_2_lut_rep_331_3_lut_4_lut (.A(stable_count[3]), .B(n21683), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21644)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2415_2_lut_rep_331_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21683), .C(stable_count[0]), 
         .D(stable_count[4]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i1_4_lut_adj_194 (.A(n21640), .B(n19937), .C(n63[2]), .D(n4), 
         .Z(stable_counting_N_2129)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_194.init = 16'h0004;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_272), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(HALL_A_OUT_c_c), .SP(clkout_c_enable_272), 
            .CK(clk_1mhz), .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(HALL_B_OUT_c_c), .SP(clkout_c_enable_272), 
            .CK(clk_1mhz), .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(HALL_C_OUT_c_c), .SP(clkout_c_enable_272), 
            .CK(clk_1mhz), .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2067[19]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2067[18]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2067[17]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2067[16]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2067[15]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2067[14]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2067[13]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2067[12]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2067[11]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2067[10]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2067[9]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2067[8]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2067[7]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2067[6]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2067[5]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2067[4]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2067[3]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2067[2]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2067[1]), .SP(clk_1mhz_enable_70), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_195 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4_adj_2426)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_195.init = 16'h7bde;
    LUT4 i2387_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2387_2_lut.init = 16'h6666;
    FD1P3AX speed__i2 (.D(speedt_19__N_2047[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2047[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2047[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2047[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2047[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2047[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2047[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2047[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2047[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2047[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2047[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2047[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2047[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2047[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2047[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2047[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2047[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2047[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2047[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i6_4_lut (.A(count[10]), .B(n12), .C(count[9]), .D(count[2]), 
         .Z(n19815)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    FD1S3IX count__i1 (.D(count_19__N_2067[1]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2067[2]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2067[3]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2067[4]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2067[5]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2067[6]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2067[7]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2067[8]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2067[9]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2067[10]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2067[11]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2067[12]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2067[13]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2067[14]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2067[15]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2067[16]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2067[17]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2067[18]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2067[19]), .CK(clk_1mhz), .CD(n4585), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    LUT4 i2401_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2401_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i5_4_lut (.A(count[3]), .B(count[8]), .C(count[13]), .D(count[0]), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i17570_4_lut (.A(n19075), .B(n20034), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_187)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17570_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_196 (.A(n19), .B(n19815), .C(n24), .D(n20), .Z(n19075)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i1_4_lut_adj_196.init = 16'hfffb;
    LUT4 i16637_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n20034)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16637_4_lut.init = 16'h7bde;
    LUT4 i6_2_lut (.A(count[17]), .B(count[12]), .Z(n19)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i11_4_lut (.A(count[5]), .B(n22), .C(n16), .D(count[16]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut (.A(count[14]), .B(count[19]), .C(count[11]), .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i9_4_lut (.A(count[15]), .B(count[18]), .C(count[1]), .D(count[4]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[6]), .B(count[7]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i2265_2_lut (.A(stable_counting), .B(stable_counting_N_2129), .Z(n4585)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2265_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_rep_369 (.A(hall3_old), .B(n4_adj_2426), .C(hall3_lat), 
         .Z(n21682)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_369.init = 16'hdede;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4_adj_2426), .C(hall3_lat), 
         .D(n63[1]), .Z(n19937)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 i2410_2_lut_rep_338_3_lut_4_lut (.A(stable_count[2]), .B(n21724), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21651)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2410_2_lut_rep_338_3_lut_4_lut.init = 16'h8000;
    LUT4 i2408_2_lut_rep_341_3_lut_4_lut (.A(stable_count[2]), .B(n21724), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21654)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2408_2_lut_rep_341_3_lut_4_lut.init = 16'h78f0;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2047[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2047[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2047[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2047[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2047[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2047[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2047[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2047[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2047[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2047[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2047[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2047[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2047[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2047[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2047[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2047[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2047[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2047[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2047[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11471), .B(n11469), .C(count_19__N_2067[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2047[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_197 (.A(n63[3]), .B(n63[6]), .C(n21644), .D(n63[2]), 
         .Z(n19814)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_197.init = 16'hfffe;
    LUT4 i16754_3_lut (.A(n21682), .B(stable_counting), .C(stable_counting_N_2129), 
         .Z(n14402)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16754_3_lut.init = 16'hc8c8;
    LUT4 i2_3_lut_rep_327_4_lut (.A(stable_count[5]), .B(n21651), .C(n63[6]), 
         .D(n63[3]), .Z(n21640)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_327_4_lut.init = 16'hfff6;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21644), .SP(stable_counting), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21654), .SP(stable_counting), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    LUT4 i2385_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2385_1_lut.init = 16'h5555;
    LUT4 i2422_3_lut_4_lut (.A(stable_count[4]), .B(n21661), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2422_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2396_2_lut_rep_370_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21683)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2396_2_lut_rep_370_3_lut.init = 16'h8080;
    FD1P3IX stable_counting_62 (.D(n22430), .SP(clk_1mhz_enable_187), .CD(n14402), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18462), 
          .S0(count_19__N_2067[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18461), .COUT(n18462), .S0(count_19__N_2067[17]), .S1(count_19__N_2067[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    LUT4 i2389_2_lut_rep_411 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21724)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2389_2_lut_rep_411.init = 16'h8888;
    LUT4 i2394_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2394_2_lut_3_lut.init = 16'h7878;
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18460), .COUT(n18461), .S0(count_19__N_2067[15]), .S1(count_19__N_2067[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18459), .COUT(n18460), .S0(count_19__N_2067[13]), .S1(count_19__N_2067[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18458), .COUT(n18459), .S0(count_19__N_2067[11]), .S1(count_19__N_2067[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18457), .COUT(n18458), .S0(count_19__N_2067[9]), .S1(count_19__N_2067[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18456), 
          .COUT(n18457), .S0(count_19__N_2067[7]), .S1(count_19__N_2067[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18455), 
          .COUT(n18456), .S0(count_19__N_2067[5]), .S1(count_19__N_2067[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18454), 
          .COUT(n18455), .S0(count_19__N_2067[3]), .S1(count_19__N_2067[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18453), 
          .COUT(n18454), .S0(count_19__N_2067[1]), .S1(count_19__N_2067[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18453), 
          .S1(count_19__N_2067[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AVG_SPEED
//

module AVG_SPEED (\speed_avg_m4[0] , clk_1mhz, \speed_m4[0] , GND_net, 
            \speed_avg_m4[1] , \speed_m4[1] , \speed_avg_m4[2] , \speed_m4[2] , 
            \speed_avg_m4[3] , \speed_m4[3] , \speed_avg_m4[4] , \speed_m4[4] , 
            \speed_avg_m4[5] , \speed_m4[5] , \speed_avg_m4[6] , \speed_m4[6] , 
            \speed_avg_m4[7] , \speed_m4[7] , \speed_avg_m4[8] , \speed_m4[8] , 
            \speed_avg_m4[9] , \speed_m4[9] , \speed_avg_m4[10] , \speed_m4[10] , 
            \speed_avg_m4[11] , \speed_m4[11] , \speed_avg_m4[12] , \speed_m4[12] , 
            \speed_avg_m4[13] , \speed_m4[13] , \speed_avg_m4[14] , \speed_m4[14] , 
            \speed_avg_m4[15] , \speed_m4[15] , \speed_avg_m4[16] , \speed_m4[16] , 
            \speed_avg_m4[17] , \speed_m4[17] , \speed_avg_m4[18] , \speed_m4[18] , 
            \speed_avg_m4[19] , \speed_m4[19] );
    output \speed_avg_m4[0] ;
    input clk_1mhz;
    input \speed_m4[0] ;
    input GND_net;
    output \speed_avg_m4[1] ;
    input \speed_m4[1] ;
    output \speed_avg_m4[2] ;
    input \speed_m4[2] ;
    output \speed_avg_m4[3] ;
    input \speed_m4[3] ;
    output \speed_avg_m4[4] ;
    input \speed_m4[4] ;
    output \speed_avg_m4[5] ;
    input \speed_m4[5] ;
    output \speed_avg_m4[6] ;
    input \speed_m4[6] ;
    output \speed_avg_m4[7] ;
    input \speed_m4[7] ;
    output \speed_avg_m4[8] ;
    input \speed_m4[8] ;
    output \speed_avg_m4[9] ;
    input \speed_m4[9] ;
    output \speed_avg_m4[10] ;
    input \speed_m4[10] ;
    output \speed_avg_m4[11] ;
    input \speed_m4[11] ;
    output \speed_avg_m4[12] ;
    input \speed_m4[12] ;
    output \speed_avg_m4[13] ;
    input \speed_m4[13] ;
    output \speed_avg_m4[14] ;
    input \speed_m4[14] ;
    output \speed_avg_m4[15] ;
    input \speed_m4[15] ;
    output \speed_avg_m4[16] ;
    input \speed_m4[16] ;
    output \speed_avg_m4[17] ;
    input \speed_m4[17] ;
    output \speed_avg_m4[18] ;
    input \speed_m4[18] ;
    output \speed_avg_m4[19] ;
    input \speed_m4[19] ;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_165;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n18542, n18541, n18540, n20166, n6;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m4[0] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2114__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_165), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114__i0.GSR = "DISABLED";
    CCU2D clk_cnt_2114_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18542), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2114_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2114_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2114_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2114_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18541), .COUT(n18542), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2114_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2114_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2114_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2114_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18540), .COUT(n18541), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2114_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2114_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2114_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2114_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18540), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2114_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2114_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2114_add_4_1.INJECT1_1 = "NO";
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m4[1] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m4[2] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m4[3] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m4[4] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m4[5] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m4[6] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m4[7] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m4[8] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m4[9] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m4[10] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m4[11] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m4[12] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m4[13] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m4[14] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m4[15] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m4[16] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m4[17] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m4[18] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m4[19] ), .SP(clk_1mhz_enable_165), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    LUT4 i17547_4_lut (.A(clk_cnt[4]), .B(n20166), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_165)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17547_4_lut.init = 16'h0004;
    LUT4 i16768_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n20166)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16768_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX clk_cnt_2114__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_165), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2114__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_165), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2114__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_165), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2114__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_165), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2114__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_165), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2114__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_165), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2114__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module SPI
//

module SPI (n22435, speed_set_m4, clkout_c, MISO_N_816, enable_m1, 
            enable_m2, enable_m3, enable_m4, clkout_c_enable_341, CS_c, 
            SCK_c, speed_set_m3, MOSI_c, GND_net, hallsense_m1, dir_m1, 
            n2872, n2908, hallsense_m2, dir_m2, n2980, n3016, clkout_c_enable_272, 
            hallsense_m3, dir_m3, n3088, n3124, rst, hallsense_m4, 
            dir_m4, n3196, n3232, n5172, speed_set_m2, speed_set_m1, 
            free_m4, n19826, free_m3, n19845, free_m2, n19830, free_m1, 
            n19843);
    input n22435;
    output [20:0]speed_set_m4;
    input clkout_c;
    output MISO_N_816;
    output enable_m1;
    output enable_m2;
    output enable_m3;
    output enable_m4;
    input clkout_c_enable_341;
    input CS_c;
    input SCK_c;
    output [20:0]speed_set_m3;
    input MOSI_c;
    input GND_net;
    input [2:0]hallsense_m1;
    input dir_m1;
    output n2872;
    output n2908;
    input [2:0]hallsense_m2;
    input dir_m2;
    output n2980;
    output n3016;
    input clkout_c_enable_272;
    input [2:0]hallsense_m3;
    input dir_m3;
    output n3088;
    output n3124;
    input rst;
    input [2:0]hallsense_m4;
    input dir_m4;
    output n3196;
    output n3232;
    output n5172;
    output [20:0]speed_set_m2;
    output [20:0]speed_set_m1;
    input free_m4;
    output n19826;
    input free_m3;
    output n19845;
    input free_m2;
    output n19830;
    input free_m1;
    output n19843;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire SCKold, CSlatched, SCKlatched, clkout_c_enable_63, clkout_c_enable_350, 
        n14152;
    wire [95:0]recv_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(68[10:21])
    wire [95:0]temp_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(70[10:21])
    wire [95:0]n193;
    
    wire MISO_N_862, n24, enable_m1_N_825, enable_m1_N_819, enable_m2_N_827, 
        enable_m3_N_834, enable_m4_N_841, CSold, n22431;
    wire [95:0]send_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(67[10:21])
    
    wire n21671, n21672;
    wire [95:0]send_buffer_95__N_442;
    
    wire MISO_N_817, n21692, n14172, MISOb, MISOb_N_852, clkout_c_enable_109, 
        n18776, n3400, n18775, n18774, n18773, n18772, n18771, 
        n18770, n18769, n21715, n21711, n18754, n3376, n18753, 
        n21704, n3496, n3472, n39, n40, n5170, n21699, n36, 
        n28, n38, n32, n18752, n18751, n18750, n18749, n18748, 
        n18747, n18746, n18745, n18744, n3448, n18743, n18742, 
        n18741, n3352, n3328, n39_adj_2394, n40_adj_2395, n36_adj_2396, 
        n28_adj_2397, n38_adj_2398, n32_adj_2399, n34, n24_adj_2400, 
        n18740, n39_adj_2401, n40_adj_2402, n36_adj_2403, n28_adj_2404, 
        n38_adj_2405, n32_adj_2406, n34_adj_2407, n24_adj_2408, n18739, 
        n18738, n18737, n3424, n39_adj_2409, n40_adj_2410, n36_adj_2411, 
        n28_adj_2412, n38_adj_2413, n32_adj_2414, n34_adj_2415, n24_adj_2416, 
        n34_adj_2417, n21690;
    wire [95:0]MISOb_N_858;
    
    wire MISOb_N_853, MISOb_N_857, n21662, n22432, n18822, n18821, 
        n18820, n18819, n18818, n18817, n18608, n18607, n18606, 
        n18605, n18816, n18604, n18815, n18814, n18603, n18602, 
        n18813, n18601, n18600, n18599, n18598, n18597, n18596, 
        n18595, n18594, n18593, n18592, n18591, n14192, n14212, 
        n18695, n18694, n18693, n18692, n18691, n18690, n18689, 
        n18688, n18794, n18793, n18792, n18791, n18790, n18789, 
        n18788, n18787, n18786, n18785;
    
    LUT4 i3_4_lut_rep_430 (.A(SCKold), .B(n22435), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_63)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut_rep_430.init = 16'h0400;
    FD1P3JX speed_set_m4_i0_i8 (.D(recv_buffer[20]), .SP(clkout_c_enable_350), 
            .PD(n14152), .CK(clkout_c), .Q(speed_set_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i8.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i0 (.D(n193[0]), .SP(clkout_c_enable_350), .CK(clkout_c), 
            .Q(temp_buffer[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i0.GSR = "DISABLED";
    FD1S3AX MISO_128 (.D(MISO_N_862), .CK(clkout_c), .Q(MISO_N_816)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISO_128.GSR = "DISABLED";
    LUT4 i3_2_lut (.A(recv_buffer[30]), .B(recv_buffer[17]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    FD1P3IX speed_set_m4_i0_i16 (.D(recv_buffer[28]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i16.GSR = "DISABLED";
    FD1P3AX enable_m1_112 (.D(enable_m1_N_819), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m1_112.GSR = "ENABLED";
    FD1P3AX enable_m2_113 (.D(enable_m2_N_827), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m2_113.GSR = "ENABLED";
    FD1P3AX enable_m3_114 (.D(enable_m3_N_834), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m3_114.GSR = "ENABLED";
    FD1P3AX enable_m4_115 (.D(enable_m4_N_841), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m4_115.GSR = "ENABLED";
    FD1P3AX CSold_116 (.D(n22431), .SP(clkout_c_enable_341), .CK(clkout_c), 
            .Q(CSold));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_116.GSR = "DISABLED";
    FD1P3AX SCKold_117 (.D(SCKlatched), .SP(clkout_c_enable_341), .CK(clkout_c), 
            .Q(SCKold));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKold_117.GSR = "DISABLED";
    FD1P3AX CSlatched_118 (.D(CS_c), .SP(clkout_c_enable_341), .CK(clkout_c), 
            .Q(CSlatched));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_118.GSR = "DISABLED";
    FD1P3AX SCKlatched_119 (.D(SCK_c), .SP(clkout_c_enable_341), .CK(clkout_c), 
            .Q(SCKlatched));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKlatched_119.GSR = "DISABLED";
    LUT4 i13132_2_lut_4_lut (.A(send_buffer[95]), .B(temp_buffer[95]), .C(n21671), 
         .D(n21672), .Z(send_buffer_95__N_442[95])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam i13132_2_lut_4_lut.init = 16'h00ca;
    FD1P3IX speed_set_m4_i0_i0 (.D(recv_buffer[12]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i0.GSR = "DISABLED";
    FD1P3AX i104_129 (.D(n21692), .SP(clkout_c_enable_341), .CK(clkout_c), 
            .Q(MISO_N_817));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i104_129.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i0 (.D(recv_buffer[33]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i0.GSR = "DISABLED";
    FD1P3AX recv_buffer_rep_5__i0 (.D(recv_buffer[1]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(n193[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer_rep_5__i0.GSR = "DISABLED";
    FD1P3AX MISOb_121 (.D(MISOb_N_852), .SP(clkout_c_enable_341), .CK(clkout_c), 
            .Q(MISOb));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISOb_121.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i17 (.D(recv_buffer[29]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i17.GSR = "DISABLED";
    FD1P3AX recv_buffer__i95 (.D(MOSI_c), .SP(clkout_c_enable_63), .CK(clkout_c), 
            .Q(recv_buffer[95])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i95.GSR = "DISABLED";
    FD1P3AX recv_buffer__i94 (.D(recv_buffer[95]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[94])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i94.GSR = "DISABLED";
    FD1P3AX recv_buffer__i93 (.D(recv_buffer[94]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i93.GSR = "DISABLED";
    FD1P3AX recv_buffer__i92 (.D(recv_buffer[93]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i92.GSR = "DISABLED";
    FD1P3AX recv_buffer__i91 (.D(recv_buffer[92]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i91.GSR = "DISABLED";
    FD1P3AX recv_buffer__i90 (.D(recv_buffer[91]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i90.GSR = "DISABLED";
    FD1P3AX recv_buffer__i89 (.D(recv_buffer[90]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i89.GSR = "DISABLED";
    FD1P3AX recv_buffer__i88 (.D(recv_buffer[89]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i88.GSR = "DISABLED";
    FD1P3AX recv_buffer__i87 (.D(recv_buffer[88]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i87.GSR = "DISABLED";
    FD1P3AX recv_buffer__i86 (.D(recv_buffer[87]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i86.GSR = "DISABLED";
    FD1P3AX recv_buffer__i85 (.D(recv_buffer[86]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i85.GSR = "DISABLED";
    FD1P3AX recv_buffer__i84 (.D(recv_buffer[85]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i84.GSR = "DISABLED";
    FD1P3AX recv_buffer__i83 (.D(recv_buffer[84]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i83.GSR = "DISABLED";
    FD1P3AX recv_buffer__i82 (.D(recv_buffer[83]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i82.GSR = "DISABLED";
    FD1P3AX recv_buffer__i81 (.D(recv_buffer[82]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i81.GSR = "DISABLED";
    FD1P3AX recv_buffer__i80 (.D(recv_buffer[81]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i80.GSR = "DISABLED";
    FD1P3AX recv_buffer__i79 (.D(recv_buffer[80]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i79.GSR = "DISABLED";
    FD1P3AX recv_buffer__i78 (.D(recv_buffer[79]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i78.GSR = "DISABLED";
    FD1P3AX recv_buffer__i77 (.D(recv_buffer[78]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i77.GSR = "DISABLED";
    FD1P3AX recv_buffer__i76 (.D(recv_buffer[77]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i76.GSR = "DISABLED";
    FD1P3AX recv_buffer__i75 (.D(recv_buffer[76]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i75.GSR = "DISABLED";
    FD1P3AX recv_buffer__i74 (.D(recv_buffer[75]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i74.GSR = "DISABLED";
    FD1P3AX recv_buffer__i73 (.D(recv_buffer[74]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i73.GSR = "DISABLED";
    FD1P3AX recv_buffer__i72 (.D(recv_buffer[73]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i72.GSR = "DISABLED";
    FD1P3AX recv_buffer__i71 (.D(recv_buffer[72]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i71.GSR = "DISABLED";
    FD1P3AX recv_buffer__i70 (.D(recv_buffer[71]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i70.GSR = "DISABLED";
    FD1P3AX recv_buffer__i69 (.D(recv_buffer[70]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i69.GSR = "DISABLED";
    FD1P3AX recv_buffer__i68 (.D(recv_buffer[69]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i68.GSR = "DISABLED";
    FD1P3AX recv_buffer__i67 (.D(recv_buffer[68]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i67.GSR = "DISABLED";
    FD1P3AX recv_buffer__i66 (.D(recv_buffer[67]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i66.GSR = "DISABLED";
    FD1P3AX recv_buffer__i65 (.D(recv_buffer[66]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i65.GSR = "DISABLED";
    FD1P3AX recv_buffer__i64 (.D(recv_buffer[65]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i64.GSR = "DISABLED";
    FD1P3AX recv_buffer__i63 (.D(recv_buffer[64]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i63.GSR = "DISABLED";
    FD1P3AX recv_buffer__i62 (.D(recv_buffer[63]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i62.GSR = "DISABLED";
    FD1P3AX recv_buffer__i61 (.D(recv_buffer[62]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i61.GSR = "DISABLED";
    FD1P3AX recv_buffer__i60 (.D(recv_buffer[61]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i60.GSR = "DISABLED";
    FD1P3AX recv_buffer__i59 (.D(recv_buffer[60]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i59.GSR = "DISABLED";
    FD1P3AX recv_buffer__i58 (.D(recv_buffer[59]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i58.GSR = "DISABLED";
    FD1P3AX recv_buffer__i57 (.D(recv_buffer[58]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i57.GSR = "DISABLED";
    FD1P3AX recv_buffer__i56 (.D(recv_buffer[57]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i56.GSR = "DISABLED";
    FD1P3AX recv_buffer__i55 (.D(recv_buffer[56]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i55.GSR = "DISABLED";
    FD1P3AX recv_buffer__i54 (.D(recv_buffer[55]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i54.GSR = "DISABLED";
    FD1P3AX recv_buffer__i53 (.D(recv_buffer[54]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i53.GSR = "DISABLED";
    FD1P3AX recv_buffer__i52 (.D(recv_buffer[53]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i52.GSR = "DISABLED";
    FD1P3AX recv_buffer__i51 (.D(recv_buffer[52]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i51.GSR = "DISABLED";
    FD1P3AX recv_buffer__i50 (.D(recv_buffer[51]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i50.GSR = "DISABLED";
    FD1P3AX recv_buffer__i49 (.D(recv_buffer[50]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i49.GSR = "DISABLED";
    FD1P3AX recv_buffer__i48 (.D(recv_buffer[49]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i48.GSR = "DISABLED";
    FD1P3AX recv_buffer__i47 (.D(recv_buffer[48]), .SP(clkout_c_enable_63), 
            .CK(clkout_c), .Q(recv_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i47.GSR = "DISABLED";
    FD1P3AX recv_buffer__i46 (.D(recv_buffer[47]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i46.GSR = "DISABLED";
    FD1P3AX recv_buffer__i45 (.D(recv_buffer[46]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i45.GSR = "DISABLED";
    FD1P3AX recv_buffer__i44 (.D(recv_buffer[45]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i44.GSR = "DISABLED";
    FD1P3AX recv_buffer__i43 (.D(recv_buffer[44]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i43.GSR = "DISABLED";
    FD1P3AX recv_buffer__i42 (.D(recv_buffer[43]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i42.GSR = "DISABLED";
    FD1P3AX recv_buffer__i41 (.D(recv_buffer[42]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i41.GSR = "DISABLED";
    FD1P3AX recv_buffer__i40 (.D(recv_buffer[41]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i40.GSR = "DISABLED";
    FD1P3AX recv_buffer__i39 (.D(recv_buffer[40]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i39.GSR = "DISABLED";
    FD1P3AX recv_buffer__i38 (.D(recv_buffer[39]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i38.GSR = "DISABLED";
    FD1P3AX recv_buffer__i37 (.D(recv_buffer[38]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i37.GSR = "DISABLED";
    FD1P3AX recv_buffer__i36 (.D(recv_buffer[37]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i36.GSR = "DISABLED";
    FD1P3AX recv_buffer__i35 (.D(recv_buffer[36]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i35.GSR = "DISABLED";
    FD1P3AX recv_buffer__i34 (.D(recv_buffer[35]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i34.GSR = "DISABLED";
    FD1P3AX recv_buffer__i33 (.D(recv_buffer[34]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i33.GSR = "DISABLED";
    FD1P3AX recv_buffer__i32 (.D(recv_buffer[33]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i32.GSR = "DISABLED";
    FD1P3AX recv_buffer__i31 (.D(recv_buffer[32]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i31.GSR = "DISABLED";
    FD1P3AX recv_buffer__i30 (.D(recv_buffer[31]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i30.GSR = "DISABLED";
    FD1P3AX recv_buffer__i29 (.D(recv_buffer[30]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i29.GSR = "DISABLED";
    FD1P3AX recv_buffer__i28 (.D(recv_buffer[29]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i28.GSR = "DISABLED";
    FD1P3AX recv_buffer__i27 (.D(recv_buffer[28]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i27.GSR = "DISABLED";
    FD1P3AX recv_buffer__i26 (.D(recv_buffer[27]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i26.GSR = "DISABLED";
    FD1P3AX recv_buffer__i25 (.D(recv_buffer[26]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i25.GSR = "DISABLED";
    FD1P3AX recv_buffer__i24 (.D(recv_buffer[25]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i24.GSR = "DISABLED";
    FD1P3AX recv_buffer__i23 (.D(recv_buffer[24]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i23.GSR = "DISABLED";
    CCU2D add_15385_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18776), 
          .S0(n3400));
    defparam add_15385_cout.INIT0 = 16'h0000;
    defparam add_15385_cout.INIT1 = 16'h0000;
    defparam add_15385_cout.INJECT1_0 = "NO";
    defparam add_15385_cout.INJECT1_1 = "NO";
    CCU2D add_15385_16 (.A0(recv_buffer[73]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[74]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18775), .COUT(n18776));
    defparam add_15385_16.INIT0 = 16'h5aaa;
    defparam add_15385_16.INIT1 = 16'h0aaa;
    defparam add_15385_16.INJECT1_0 = "NO";
    defparam add_15385_16.INJECT1_1 = "NO";
    FD1P3AX recv_buffer__i22 (.D(recv_buffer[23]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i22.GSR = "DISABLED";
    FD1P3AX recv_buffer__i21 (.D(recv_buffer[22]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i21.GSR = "DISABLED";
    FD1P3AX recv_buffer__i20 (.D(recv_buffer[21]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i20.GSR = "DISABLED";
    FD1P3AX recv_buffer__i19 (.D(recv_buffer[20]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i19.GSR = "DISABLED";
    FD1P3AX recv_buffer__i18 (.D(recv_buffer[19]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i18.GSR = "DISABLED";
    FD1P3AX recv_buffer__i17 (.D(recv_buffer[18]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i17.GSR = "DISABLED";
    FD1P3AX recv_buffer__i16 (.D(recv_buffer[17]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i16.GSR = "DISABLED";
    FD1P3AX recv_buffer__i15 (.D(recv_buffer[16]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i15.GSR = "DISABLED";
    FD1P3AX recv_buffer__i14 (.D(recv_buffer[15]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i14.GSR = "DISABLED";
    FD1P3AX recv_buffer__i13 (.D(recv_buffer[14]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i13.GSR = "DISABLED";
    FD1P3AX recv_buffer__i12 (.D(recv_buffer[13]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i12.GSR = "DISABLED";
    FD1P3AX recv_buffer__i11 (.D(recv_buffer[12]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i11.GSR = "DISABLED";
    FD1P3AX recv_buffer__i10 (.D(recv_buffer[11]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i10.GSR = "DISABLED";
    FD1P3AX recv_buffer__i9 (.D(recv_buffer[10]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i9.GSR = "DISABLED";
    FD1P3AX recv_buffer__i8 (.D(recv_buffer[9]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i8.GSR = "DISABLED";
    FD1P3AX recv_buffer__i7 (.D(recv_buffer[8]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i7.GSR = "DISABLED";
    FD1P3AX recv_buffer__i6 (.D(recv_buffer[7]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i6.GSR = "DISABLED";
    FD1P3AX recv_buffer__i5 (.D(recv_buffer[6]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i5.GSR = "DISABLED";
    FD1P3AX recv_buffer__i4 (.D(recv_buffer[5]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i4.GSR = "DISABLED";
    FD1P3AX recv_buffer__i3 (.D(recv_buffer[4]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i3.GSR = "DISABLED";
    FD1P3AX recv_buffer__i2 (.D(recv_buffer[3]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i2.GSR = "DISABLED";
    FD1P3AX recv_buffer__i1 (.D(recv_buffer[2]), .SP(clkout_c_enable_109), 
            .CK(clkout_c), .Q(recv_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i1.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i95 (.D(recv_buffer[95]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[95])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i95.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i94 (.D(recv_buffer[94]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[94])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i94.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i93 (.D(recv_buffer[93]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i93.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i92 (.D(recv_buffer[92]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i92.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i91 (.D(recv_buffer[91]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i91.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i90 (.D(recv_buffer[90]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i90.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i89 (.D(recv_buffer[89]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i89.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i88 (.D(recv_buffer[88]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i88.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i87 (.D(recv_buffer[87]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i87.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i86 (.D(recv_buffer[86]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i86.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i85 (.D(recv_buffer[85]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i85.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i84 (.D(recv_buffer[84]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i84.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i83 (.D(recv_buffer[83]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i83.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i82 (.D(recv_buffer[82]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i82.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i81 (.D(recv_buffer[81]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i81.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i80 (.D(recv_buffer[80]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i80.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i79 (.D(recv_buffer[79]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i79.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i78 (.D(recv_buffer[78]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i78.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i77 (.D(recv_buffer[77]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i77.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i76 (.D(recv_buffer[76]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i76.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i75 (.D(recv_buffer[75]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i75.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i74 (.D(recv_buffer[74]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i74.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i73 (.D(recv_buffer[73]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i73.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i72 (.D(recv_buffer[72]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i72.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i71 (.D(recv_buffer[71]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i71.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i70 (.D(recv_buffer[70]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i70.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i69 (.D(recv_buffer[69]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i69.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i68 (.D(recv_buffer[68]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i68.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i67 (.D(recv_buffer[67]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i67.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i66 (.D(recv_buffer[66]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i66.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i65 (.D(recv_buffer[65]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i65.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i64 (.D(recv_buffer[64]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i64.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i63 (.D(recv_buffer[63]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i63.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i62 (.D(recv_buffer[62]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i62.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i61 (.D(recv_buffer[61]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i61.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i60 (.D(recv_buffer[60]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i60.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i59 (.D(recv_buffer[59]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i59.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i58 (.D(recv_buffer[58]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i58.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i57 (.D(recv_buffer[57]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i57.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i56 (.D(recv_buffer[56]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i56.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i55 (.D(recv_buffer[55]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i55.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i54 (.D(recv_buffer[54]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i54.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i53 (.D(recv_buffer[53]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i53.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i52 (.D(recv_buffer[52]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i52.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i51 (.D(recv_buffer[51]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i51.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i50 (.D(recv_buffer[50]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i50.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i49 (.D(recv_buffer[49]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i49.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i48 (.D(recv_buffer[48]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i48.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i47 (.D(recv_buffer[47]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i47.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i46 (.D(recv_buffer[46]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i46.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i45 (.D(recv_buffer[45]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i45.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i44 (.D(recv_buffer[44]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i44.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i43 (.D(recv_buffer[43]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i43.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i42 (.D(recv_buffer[42]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i42.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i41 (.D(recv_buffer[41]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i41.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i40 (.D(recv_buffer[40]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i40.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i39 (.D(recv_buffer[39]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i39.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i38 (.D(recv_buffer[38]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i38.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i37 (.D(recv_buffer[37]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i37.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i36 (.D(recv_buffer[36]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i36.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i35 (.D(recv_buffer[35]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i35.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i34 (.D(recv_buffer[34]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i34.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i33 (.D(recv_buffer[33]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i33.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i32 (.D(recv_buffer[32]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i32.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i31 (.D(recv_buffer[31]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i31.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i30 (.D(recv_buffer[30]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i30.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i29 (.D(recv_buffer[29]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i29.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i28 (.D(recv_buffer[28]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i28.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i27 (.D(recv_buffer[27]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i27.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i26 (.D(recv_buffer[26]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i26.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i25 (.D(recv_buffer[25]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i25.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i24 (.D(recv_buffer[24]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i24.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i23 (.D(recv_buffer[23]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i23.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i22 (.D(recv_buffer[22]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i22.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i21 (.D(recv_buffer[21]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i21.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i20 (.D(recv_buffer[20]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i20.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i19 (.D(recv_buffer[19]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i19.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i18 (.D(recv_buffer[18]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i18.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i17 (.D(recv_buffer[17]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i17.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i16 (.D(recv_buffer[16]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i16.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i15 (.D(recv_buffer[15]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i15.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i14 (.D(recv_buffer[14]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i14.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i13 (.D(recv_buffer[13]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i13.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i12 (.D(recv_buffer[12]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i12.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i11 (.D(recv_buffer[11]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i11.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i10 (.D(recv_buffer[10]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i10.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i9 (.D(recv_buffer[9]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i9.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i8 (.D(recv_buffer[8]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i8.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i7 (.D(recv_buffer[7]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i6 (.D(recv_buffer[6]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i5 (.D(recv_buffer[5]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i5.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i4 (.D(recv_buffer[4]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i4.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i3 (.D(recv_buffer[3]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i2 (.D(recv_buffer[2]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i1 (.D(recv_buffer[1]), .SP(clkout_c_enable_350), 
            .CK(clkout_c), .Q(temp_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i1.GSR = "DISABLED";
    CCU2D add_15385_14 (.A0(recv_buffer[71]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[72]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18774), .COUT(n18775));
    defparam add_15385_14.INIT0 = 16'h5aaa;
    defparam add_15385_14.INIT1 = 16'h5aaa;
    defparam add_15385_14.INJECT1_0 = "NO";
    defparam add_15385_14.INJECT1_1 = "NO";
    CCU2D add_15385_12 (.A0(recv_buffer[69]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[70]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18773), .COUT(n18774));
    defparam add_15385_12.INIT0 = 16'h5aaa;
    defparam add_15385_12.INIT1 = 16'h5aaa;
    defparam add_15385_12.INJECT1_0 = "NO";
    defparam add_15385_12.INJECT1_1 = "NO";
    CCU2D add_15385_10 (.A0(recv_buffer[67]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[68]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18772), .COUT(n18773));
    defparam add_15385_10.INIT0 = 16'h5555;
    defparam add_15385_10.INIT1 = 16'h5aaa;
    defparam add_15385_10.INJECT1_0 = "NO";
    defparam add_15385_10.INJECT1_1 = "NO";
    CCU2D add_15385_8 (.A0(recv_buffer[65]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[66]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18771), .COUT(n18772));
    defparam add_15385_8.INIT0 = 16'h5aaa;
    defparam add_15385_8.INIT1 = 16'h5aaa;
    defparam add_15385_8.INJECT1_0 = "NO";
    defparam add_15385_8.INJECT1_1 = "NO";
    CCU2D add_15385_6 (.A0(recv_buffer[63]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[64]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18770), .COUT(n18771));
    defparam add_15385_6.INIT0 = 16'h5555;
    defparam add_15385_6.INIT1 = 16'h5555;
    defparam add_15385_6.INJECT1_0 = "NO";
    defparam add_15385_6.INJECT1_1 = "NO";
    CCU2D add_15385_4 (.A0(recv_buffer[61]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[62]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18769), .COUT(n18770));
    defparam add_15385_4.INIT0 = 16'h5aaa;
    defparam add_15385_4.INIT1 = 16'h5555;
    defparam add_15385_4.INJECT1_0 = "NO";
    defparam add_15385_4.INJECT1_1 = "NO";
    CCU2D add_15385_2 (.A0(recv_buffer[59]), .B0(recv_buffer[58]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[60]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18769));
    defparam add_15385_2.INIT0 = 16'h7000;
    defparam add_15385_2.INIT1 = 16'h5aaa;
    defparam add_15385_2.INJECT1_0 = "NO";
    defparam add_15385_2.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(hallsense_m1[2]), .B(n21715), .C(dir_m1), .D(hallsense_m1[1]), 
         .Z(n2872)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut.init = 16'h4008;
    LUT4 i1_4_lut_adj_160 (.A(hallsense_m1[1]), .B(n21715), .C(dir_m1), 
         .D(hallsense_m1[0]), .Z(n2908)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_160.init = 16'h4008;
    LUT4 i1_4_lut_adj_161 (.A(hallsense_m2[2]), .B(n21711), .C(dir_m2), 
         .D(hallsense_m2[1]), .Z(n2980)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_161.init = 16'h4008;
    LUT4 i1_4_lut_adj_162 (.A(hallsense_m2[1]), .B(n21711), .C(dir_m2), 
         .D(hallsense_m2[0]), .Z(n3016)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_162.init = 16'h4008;
    CCU2D add_15386_21 (.A0(recv_buffer[74]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18754), .S1(n3376));
    defparam add_15386_21.INIT0 = 16'h5555;
    defparam add_15386_21.INIT1 = 16'h0000;
    defparam add_15386_21.INJECT1_0 = "NO";
    defparam add_15386_21.INJECT1_1 = "NO";
    CCU2D add_15386_19 (.A0(recv_buffer[72]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[73]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18753), .COUT(n18754));
    defparam add_15386_19.INIT0 = 16'hf555;
    defparam add_15386_19.INIT1 = 16'hf555;
    defparam add_15386_19.INJECT1_0 = "NO";
    defparam add_15386_19.INJECT1_1 = "NO";
    FD1P3AX send_buffer_i0_i1 (.D(send_buffer_95__N_442[1]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_163 (.A(hallsense_m3[2]), .B(n21704), .C(dir_m3), 
         .D(hallsense_m3[1]), .Z(n3088)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_163.init = 16'h4008;
    LUT4 i1_4_lut_adj_164 (.A(hallsense_m3[1]), .B(n21704), .C(dir_m3), 
         .D(hallsense_m3[0]), .Z(n3124)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_164.init = 16'h4008;
    LUT4 i2_4_lut (.A(n3496), .B(n3472), .C(n39), .D(n40), .Z(enable_m4_N_841)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    FD1P3AX send_buffer_i0_i2 (.D(send_buffer_95__N_442[2]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i3 (.D(send_buffer_95__N_442[3]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i4 (.D(send_buffer_95__N_442[4]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i4.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i5 (.D(send_buffer_95__N_442[5]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i5.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i6 (.D(send_buffer_95__N_442[6]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i7 (.D(send_buffer_95__N_442[7]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i8 (.D(send_buffer_95__N_442[8]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i8.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i9 (.D(send_buffer_95__N_442[9]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i9.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i10 (.D(send_buffer_95__N_442[10]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i10.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i11 (.D(send_buffer_95__N_442[11]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i11.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i12 (.D(send_buffer_95__N_442[12]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i12.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i13 (.D(send_buffer_95__N_442[13]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i13.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i14 (.D(send_buffer_95__N_442[14]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i14.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i15 (.D(send_buffer_95__N_442[15]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i15.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i16 (.D(send_buffer_95__N_442[16]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i16.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i17 (.D(send_buffer_95__N_442[17]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i17.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i18 (.D(send_buffer_95__N_442[18]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i18.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i19 (.D(send_buffer_95__N_442[19]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i19.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i20 (.D(send_buffer_95__N_442[20]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i20.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i21 (.D(send_buffer_95__N_442[21]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i21.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i22 (.D(send_buffer_95__N_442[22]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i22.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i23 (.D(send_buffer_95__N_442[23]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i23.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i24 (.D(send_buffer_95__N_442[24]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i24.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i25 (.D(send_buffer_95__N_442[25]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i25.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i26 (.D(send_buffer_95__N_442[26]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i26.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i27 (.D(send_buffer_95__N_442[27]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i27.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i28 (.D(send_buffer_95__N_442[28]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i28.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i29 (.D(send_buffer_95__N_442[29]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i29.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i30 (.D(send_buffer_95__N_442[30]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i30.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i31 (.D(send_buffer_95__N_442[31]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i31.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i32 (.D(send_buffer_95__N_442[32]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i32.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i33 (.D(send_buffer_95__N_442[33]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i33.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i34 (.D(send_buffer_95__N_442[34]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i34.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i35 (.D(send_buffer_95__N_442[35]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i35.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i36 (.D(send_buffer_95__N_442[36]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i36.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i37 (.D(send_buffer_95__N_442[37]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i37.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i38 (.D(send_buffer_95__N_442[38]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i38.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i39 (.D(send_buffer_95__N_442[39]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i39.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i40 (.D(send_buffer_95__N_442[40]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i40.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i41 (.D(send_buffer_95__N_442[41]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i41.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i42 (.D(send_buffer_95__N_442[42]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i42.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i43 (.D(send_buffer_95__N_442[43]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i43.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i44 (.D(send_buffer_95__N_442[44]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i44.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i45 (.D(send_buffer_95__N_442[45]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i45.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i46 (.D(send_buffer_95__N_442[46]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i46.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i47 (.D(send_buffer_95__N_442[47]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i47.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i48 (.D(send_buffer_95__N_442[48]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i48.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i49 (.D(send_buffer_95__N_442[49]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i49.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i50 (.D(send_buffer_95__N_442[50]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i50.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i51 (.D(send_buffer_95__N_442[51]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i51.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i52 (.D(send_buffer_95__N_442[52]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i52.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i53 (.D(send_buffer_95__N_442[53]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i53.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i54 (.D(send_buffer_95__N_442[54]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i54.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i55 (.D(send_buffer_95__N_442[55]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i55.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i56 (.D(send_buffer_95__N_442[56]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i56.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i57 (.D(send_buffer_95__N_442[57]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i57.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i58 (.D(send_buffer_95__N_442[58]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i58.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i59 (.D(send_buffer_95__N_442[59]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i59.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i60 (.D(send_buffer_95__N_442[60]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i60.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i61 (.D(send_buffer_95__N_442[61]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i61.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i62 (.D(send_buffer_95__N_442[62]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i62.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i63 (.D(send_buffer_95__N_442[63]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i63.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i64 (.D(send_buffer_95__N_442[64]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i64.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i65 (.D(send_buffer_95__N_442[65]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i65.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i66 (.D(send_buffer_95__N_442[66]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i66.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i67 (.D(send_buffer_95__N_442[67]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i67.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i68 (.D(send_buffer_95__N_442[68]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i68.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i69 (.D(send_buffer_95__N_442[69]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i69.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i70 (.D(send_buffer_95__N_442[70]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i70.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i71 (.D(send_buffer_95__N_442[71]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i71.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i72 (.D(send_buffer_95__N_442[72]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i72.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i73 (.D(send_buffer_95__N_442[73]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i73.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i74 (.D(send_buffer_95__N_442[74]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i74.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i75 (.D(send_buffer_95__N_442[75]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i75.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i76 (.D(send_buffer_95__N_442[76]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i76.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i77 (.D(send_buffer_95__N_442[77]), .SP(clkout_c_enable_272), 
            .CK(clkout_c), .Q(send_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i77.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i78 (.D(send_buffer_95__N_442[78]), .SP(clkout_c_enable_341), 
            .CK(clkout_c), .Q(send_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i78.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i79 (.D(send_buffer_95__N_442[79]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i79.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i80 (.D(send_buffer_95__N_442[80]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i80.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i81 (.D(send_buffer_95__N_442[81]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i81.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i82 (.D(send_buffer_95__N_442[82]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i82.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i83 (.D(send_buffer_95__N_442[83]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i83.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i84 (.D(send_buffer_95__N_442[84]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i84.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i85 (.D(send_buffer_95__N_442[85]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i85.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i86 (.D(send_buffer_95__N_442[86]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i86.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i87 (.D(send_buffer_95__N_442[87]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i87.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i88 (.D(send_buffer_95__N_442[88]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i88.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i89 (.D(send_buffer_95__N_442[89]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i89.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i90 (.D(send_buffer_95__N_442[90]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i90.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i91 (.D(send_buffer_95__N_442[91]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i91.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i92 (.D(send_buffer_95__N_442[92]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i92.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i93 (.D(send_buffer_95__N_442[93]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i93.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i94 (.D(send_buffer_95__N_442[94]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[94])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i94.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i95 (.D(send_buffer_95__N_442[95]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[95])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i95.GSR = "DISABLED";
    LUT4 i2744_2_lut (.A(MISO_N_816), .B(MISO_N_817), .Z(n5170)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    defparam i2744_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_165 (.A(hallsense_m4[2]), .B(n21699), .C(dir_m4), 
         .D(hallsense_m4[1]), .Z(n3196)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_165.init = 16'h4008;
    LUT4 i18_4_lut (.A(recv_buffer[25]), .B(n36), .C(n28), .D(recv_buffer[24]), 
         .Z(n39)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(recv_buffer[27]), .B(n38), .C(n32), .D(recv_buffer[22]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_166 (.A(hallsense_m4[1]), .B(n21699), .C(dir_m4), 
         .D(hallsense_m4[0]), .Z(n3232)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_166.init = 16'h4008;
    CCU2D add_15386_17 (.A0(recv_buffer[70]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[71]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18752), .COUT(n18753));
    defparam add_15386_17.INIT0 = 16'hf555;
    defparam add_15386_17.INIT1 = 16'hf555;
    defparam add_15386_17.INJECT1_0 = "NO";
    defparam add_15386_17.INJECT1_1 = "NO";
    CCU2D add_15386_15 (.A0(recv_buffer[68]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[69]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18751), .COUT(n18752));
    defparam add_15386_15.INIT0 = 16'hf555;
    defparam add_15386_15.INIT1 = 16'hf555;
    defparam add_15386_15.INJECT1_0 = "NO";
    defparam add_15386_15.INJECT1_1 = "NO";
    CCU2D add_15386_13 (.A0(recv_buffer[66]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[67]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18750), .COUT(n18751));
    defparam add_15386_13.INIT0 = 16'hf555;
    defparam add_15386_13.INIT1 = 16'h0aaa;
    defparam add_15386_13.INJECT1_0 = "NO";
    defparam add_15386_13.INJECT1_1 = "NO";
    CCU2D add_15386_11 (.A0(recv_buffer[64]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[65]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18749), .COUT(n18750));
    defparam add_15386_11.INIT0 = 16'h0aaa;
    defparam add_15386_11.INIT1 = 16'hf555;
    defparam add_15386_11.INJECT1_0 = "NO";
    defparam add_15386_11.INJECT1_1 = "NO";
    CCU2D add_15386_9 (.A0(recv_buffer[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18748), .COUT(n18749));
    defparam add_15386_9.INIT0 = 16'h0aaa;
    defparam add_15386_9.INIT1 = 16'h0aaa;
    defparam add_15386_9.INJECT1_0 = "NO";
    defparam add_15386_9.INJECT1_1 = "NO";
    CCU2D add_15386_7 (.A0(recv_buffer[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18747), .COUT(n18748));
    defparam add_15386_7.INIT0 = 16'hf555;
    defparam add_15386_7.INIT1 = 16'hf555;
    defparam add_15386_7.INJECT1_0 = "NO";
    defparam add_15386_7.INJECT1_1 = "NO";
    CCU2D add_15386_5 (.A0(recv_buffer[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18746), .COUT(n18747));
    defparam add_15386_5.INIT0 = 16'h0aaa;
    defparam add_15386_5.INIT1 = 16'hf555;
    defparam add_15386_5.INJECT1_0 = "NO";
    defparam add_15386_5.INJECT1_1 = "NO";
    CCU2D add_15386_3 (.A0(recv_buffer[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18745), .COUT(n18746));
    defparam add_15386_3.INIT0 = 16'hf555;
    defparam add_15386_3.INIT1 = 16'hf555;
    defparam add_15386_3.INJECT1_0 = "NO";
    defparam add_15386_3.INJECT1_1 = "NO";
    CCU2D add_15386_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[54]), .B1(recv_buffer[55]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18745));
    defparam add_15386_1.INIT0 = 16'hF000;
    defparam add_15386_1.INIT1 = 16'ha666;
    defparam add_15386_1.INJECT1_0 = "NO";
    defparam add_15386_1.INJECT1_1 = "NO";
    CCU2D add_15387_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18744), 
          .S0(n3448));
    defparam add_15387_cout.INIT0 = 16'h0000;
    defparam add_15387_cout.INIT1 = 16'h0000;
    defparam add_15387_cout.INJECT1_0 = "NO";
    defparam add_15387_cout.INJECT1_1 = "NO";
    CCU2D add_15387_16 (.A0(recv_buffer[52]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[53]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18743), .COUT(n18744));
    defparam add_15387_16.INIT0 = 16'h5aaa;
    defparam add_15387_16.INIT1 = 16'h0aaa;
    defparam add_15387_16.INJECT1_0 = "NO";
    defparam add_15387_16.INJECT1_1 = "NO";
    CCU2D add_15387_14 (.A0(recv_buffer[50]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[51]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18742), .COUT(n18743));
    defparam add_15387_14.INIT0 = 16'h5aaa;
    defparam add_15387_14.INIT1 = 16'h5aaa;
    defparam add_15387_14.INJECT1_0 = "NO";
    defparam add_15387_14.INJECT1_1 = "NO";
    LUT4 CSold_I_0_136_2_lut (.A(CSold), .B(CSlatched), .Z(enable_m1_N_825)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam CSold_I_0_136_2_lut.init = 16'h8888;
    CCU2D add_15387_12 (.A0(recv_buffer[48]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[49]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18741), .COUT(n18742));
    defparam add_15387_12.INIT0 = 16'h5aaa;
    defparam add_15387_12.INIT1 = 16'h5aaa;
    defparam add_15387_12.INJECT1_0 = "NO";
    defparam add_15387_12.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_167 (.A(n3352), .B(n3328), .C(n39_adj_2394), .D(n40_adj_2395), 
         .Z(enable_m1_N_819)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_167.init = 16'h8880;
    LUT4 i18_4_lut_adj_168 (.A(recv_buffer[88]), .B(n36_adj_2396), .C(n28_adj_2397), 
         .D(recv_buffer[87]), .Z(n39_adj_2394)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_168.init = 16'hfffe;
    LUT4 i19_4_lut_adj_169 (.A(recv_buffer[90]), .B(n38_adj_2398), .C(n32_adj_2399), 
         .D(recv_buffer[85]), .Z(n40_adj_2395)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_169.init = 16'hfffe;
    LUT4 i15_4_lut (.A(recv_buffer[75]), .B(recv_buffer[82]), .C(recv_buffer[92]), 
         .D(recv_buffer[86]), .Z(n36_adj_2396)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(recv_buffer[76]), .B(recv_buffer[77]), .Z(n28_adj_2397)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(recv_buffer[83]), .B(n34), .C(n24_adj_2400), .D(recv_buffer[91]), 
         .Z(n38_adj_2398)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    CCU2D add_15387_10 (.A0(recv_buffer[46]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[47]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18740), .COUT(n18741));
    defparam add_15387_10.INIT0 = 16'h5555;
    defparam add_15387_10.INIT1 = 16'h5aaa;
    defparam add_15387_10.INJECT1_0 = "NO";
    defparam add_15387_10.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(recv_buffer[81]), .B(recv_buffer[78]), .C(recv_buffer[89]), 
         .Z(n32_adj_2399)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(recv_buffer[95]), .B(recv_buffer[94]), .C(recv_buffer[84]), 
         .D(recv_buffer[79]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut_adj_170 (.A(recv_buffer[93]), .B(recv_buffer[80]), .Z(n24_adj_2400)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_170.init = 16'heeee;
    LUT4 i2_4_lut_adj_171 (.A(n3400), .B(n3376), .C(n39_adj_2401), .D(n40_adj_2402), 
         .Z(enable_m2_N_827)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_171.init = 16'h8880;
    LUT4 i18_4_lut_adj_172 (.A(recv_buffer[67]), .B(n36_adj_2403), .C(n28_adj_2404), 
         .D(recv_buffer[66]), .Z(n39_adj_2401)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_172.init = 16'hfffe;
    LUT4 i19_4_lut_adj_173 (.A(recv_buffer[69]), .B(n38_adj_2405), .C(n32_adj_2406), 
         .D(recv_buffer[64]), .Z(n40_adj_2402)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_173.init = 16'hfffe;
    LUT4 i15_4_lut_adj_174 (.A(recv_buffer[54]), .B(recv_buffer[61]), .C(recv_buffer[71]), 
         .D(recv_buffer[65]), .Z(n36_adj_2403)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_174.init = 16'hfffe;
    LUT4 i7_2_lut_adj_175 (.A(recv_buffer[55]), .B(recv_buffer[56]), .Z(n28_adj_2404)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_175.init = 16'heeee;
    LUT4 i17_4_lut_adj_176 (.A(recv_buffer[62]), .B(n34_adj_2407), .C(n24_adj_2408), 
         .D(recv_buffer[70]), .Z(n38_adj_2405)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_176.init = 16'hfffe;
    LUT4 i11_3_lut_adj_177 (.A(recv_buffer[60]), .B(recv_buffer[57]), .C(recv_buffer[68]), 
         .Z(n32_adj_2406)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_177.init = 16'hfefe;
    LUT4 i13_4_lut_adj_178 (.A(recv_buffer[74]), .B(recv_buffer[73]), .C(recv_buffer[63]), 
         .D(recv_buffer[58]), .Z(n34_adj_2407)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_178.init = 16'hfffe;
    CCU2D add_15387_8 (.A0(recv_buffer[44]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[45]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18739), .COUT(n18740));
    defparam add_15387_8.INIT0 = 16'h5aaa;
    defparam add_15387_8.INIT1 = 16'h5aaa;
    defparam add_15387_8.INJECT1_0 = "NO";
    defparam add_15387_8.INJECT1_1 = "NO";
    CCU2D add_15387_6 (.A0(recv_buffer[42]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[43]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18738), .COUT(n18739));
    defparam add_15387_6.INIT0 = 16'h5555;
    defparam add_15387_6.INIT1 = 16'h5555;
    defparam add_15387_6.INJECT1_0 = "NO";
    defparam add_15387_6.INJECT1_1 = "NO";
    LUT4 i3_2_lut_adj_179 (.A(recv_buffer[72]), .B(recv_buffer[59]), .Z(n24_adj_2408)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_179.init = 16'heeee;
    CCU2D add_15387_4 (.A0(recv_buffer[40]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[41]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18737), .COUT(n18738));
    defparam add_15387_4.INIT0 = 16'h5aaa;
    defparam add_15387_4.INIT1 = 16'h5555;
    defparam add_15387_4.INJECT1_0 = "NO";
    defparam add_15387_4.INJECT1_1 = "NO";
    CCU2D add_15387_2 (.A0(recv_buffer[38]), .B0(recv_buffer[37]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[39]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18737));
    defparam add_15387_2.INIT0 = 16'h7000;
    defparam add_15387_2.INIT1 = 16'h5aaa;
    defparam add_15387_2.INJECT1_0 = "NO";
    defparam add_15387_2.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_180 (.A(n3448), .B(n3424), .C(n39_adj_2409), .D(n40_adj_2410), 
         .Z(enable_m3_N_834)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_180.init = 16'h8880;
    LUT4 i18_4_lut_adj_181 (.A(recv_buffer[46]), .B(n36_adj_2411), .C(n28_adj_2412), 
         .D(recv_buffer[45]), .Z(n39_adj_2409)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_181.init = 16'hfffe;
    LUT4 i19_4_lut_adj_182 (.A(recv_buffer[48]), .B(n38_adj_2413), .C(n32_adj_2414), 
         .D(recv_buffer[43]), .Z(n40_adj_2410)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_182.init = 16'hfffe;
    LUT4 i15_4_lut_adj_183 (.A(recv_buffer[33]), .B(recv_buffer[40]), .C(recv_buffer[50]), 
         .D(recv_buffer[44]), .Z(n36_adj_2411)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_183.init = 16'hfffe;
    LUT4 i7_2_lut_adj_184 (.A(recv_buffer[34]), .B(recv_buffer[35]), .Z(n28_adj_2412)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_184.init = 16'heeee;
    LUT4 i17_4_lut_adj_185 (.A(recv_buffer[41]), .B(n34_adj_2415), .C(n24_adj_2416), 
         .D(recv_buffer[49]), .Z(n38_adj_2413)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_185.init = 16'hfffe;
    LUT4 i11_3_lut_adj_186 (.A(recv_buffer[39]), .B(recv_buffer[36]), .C(recv_buffer[47]), 
         .Z(n32_adj_2414)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_186.init = 16'hfefe;
    LUT4 i13_4_lut_adj_187 (.A(recv_buffer[53]), .B(recv_buffer[52]), .C(recv_buffer[42]), 
         .D(recv_buffer[37]), .Z(n34_adj_2415)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_187.init = 16'hfffe;
    LUT4 i3_2_lut_adj_188 (.A(recv_buffer[51]), .B(recv_buffer[38]), .Z(n24_adj_2416)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_188.init = 16'heeee;
    LUT4 i3_4_lut (.A(SCKold), .B(n22435), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_109)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i15_4_lut_adj_189 (.A(recv_buffer[12]), .B(recv_buffer[19]), .C(recv_buffer[29]), 
         .D(recv_buffer[23]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_189.init = 16'hfffe;
    LUT4 i7_2_lut_adj_190 (.A(recv_buffer[13]), .B(recv_buffer[14]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_190.init = 16'heeee;
    LUT4 i17_4_lut_adj_191 (.A(recv_buffer[20]), .B(n34_adj_2417), .C(n24), 
         .D(recv_buffer[28]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_191.init = 16'hfffe;
    LUT4 SCKold_I_0_2_lut_rep_377 (.A(SCKold), .B(SCKlatched), .Z(n21690)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(193[8:45])
    defparam SCKold_I_0_2_lut_rep_377.init = 16'h2222;
    LUT4 MISOb_N_853_I_0_3_lut_4_lut (.A(SCKold), .B(SCKlatched), .C(MISOb_N_858[1]), 
         .D(MISOb_N_853), .Z(MISOb_N_857)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(193[8:45])
    defparam MISOb_N_853_I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11_3_lut_adj_192 (.A(recv_buffer[18]), .B(recv_buffer[15]), .C(recv_buffer[26]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_192.init = 16'hfefe;
    LUT4 CSlatched_I_0_1_lut_rep_379 (.A(CSlatched), .Z(n21692)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam CSlatched_I_0_1_lut_rep_379.init = 16'h5555;
    LUT4 mux_9_i96_3_lut_rep_349_4_lut_4_lut (.A(n22431), .B(send_buffer[95]), 
         .C(temp_buffer[95]), .D(CSold), .Z(n21662)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i96_3_lut_rep_349_4_lut_4_lut.init = 16'hd8cc;
    LUT4 CSold_I_0_2_lut_rep_358_2_lut (.A(n22431), .B(n22432), .Z(n21671)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam CSold_I_0_2_lut_rep_358_2_lut.init = 16'h4444;
    LUT4 i2743_1_lut (.A(MISO_N_817), .Z(n5172)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    defparam i2743_1_lut.init = 16'h5555;
    LUT4 MISOb_I_0_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb), .C(temp_buffer[0]), 
         .D(n22432), .Z(MISOb_N_853)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam MISOb_I_0_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i2_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[1]), .C(temp_buffer[1]), 
         .D(n22432), .Z(MISOb_N_858[1])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i2_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i3_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[2]), .C(temp_buffer[2]), 
         .D(n22432), .Z(MISOb_N_858[2])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i3_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i4_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[3]), .C(temp_buffer[3]), 
         .D(n22432), .Z(MISOb_N_858[3])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i4_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i5_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[4]), .C(temp_buffer[4]), 
         .D(n22432), .Z(MISOb_N_858[4])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i5_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i6_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[5]), .C(temp_buffer[5]), 
         .D(n22432), .Z(MISOb_N_858[5])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i6_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i7_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[6]), .C(temp_buffer[6]), 
         .D(n22432), .Z(MISOb_N_858[6])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i7_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i8_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[7]), .C(temp_buffer[7]), 
         .D(n22432), .Z(MISOb_N_858[7])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i8_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i9_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[8]), .C(temp_buffer[8]), 
         .D(n22432), .Z(MISOb_N_858[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i10_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[9]), .C(temp_buffer[9]), 
         .D(n22432), .Z(MISOb_N_858[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i11_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[10]), .C(temp_buffer[10]), 
         .D(n22432), .Z(MISOb_N_858[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i12_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[11]), .C(temp_buffer[11]), 
         .D(n22432), .Z(MISOb_N_858[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i13_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[12]), .C(temp_buffer[12]), 
         .D(n22432), .Z(MISOb_N_858[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i14_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[13]), .C(temp_buffer[13]), 
         .D(n22432), .Z(MISOb_N_858[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i15_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[14]), .C(temp_buffer[14]), 
         .D(n22432), .Z(MISOb_N_858[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i16_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[15]), .C(temp_buffer[15]), 
         .D(n22432), .Z(MISOb_N_858[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i17_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[16]), .C(temp_buffer[16]), 
         .D(n22432), .Z(MISOb_N_858[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i18_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[17]), .C(temp_buffer[17]), 
         .D(n22432), .Z(MISOb_N_858[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i19_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[18]), .C(temp_buffer[18]), 
         .D(n22432), .Z(MISOb_N_858[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i20_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[19]), .C(temp_buffer[19]), 
         .D(n22432), .Z(MISOb_N_858[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_21 (.A0(recv_buffer[95]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18822), .S1(n3328));
    defparam add_15368_21.INIT0 = 16'h5555;
    defparam add_15368_21.INIT1 = 16'h0000;
    defparam add_15368_21.INJECT1_0 = "NO";
    defparam add_15368_21.INJECT1_1 = "NO";
    LUT4 mux_9_i21_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[20]), .C(temp_buffer[20]), 
         .D(n22432), .Z(MISOb_N_858[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i22_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[21]), .C(temp_buffer[21]), 
         .D(n22432), .Z(MISOb_N_858[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i23_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[22]), .C(temp_buffer[22]), 
         .D(n22432), .Z(MISOb_N_858[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i24_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[23]), .C(temp_buffer[23]), 
         .D(n22432), .Z(MISOb_N_858[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i25_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[24]), .C(temp_buffer[24]), 
         .D(n22432), .Z(MISOb_N_858[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i26_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[25]), .C(temp_buffer[25]), 
         .D(n22432), .Z(MISOb_N_858[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i27_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[26]), .C(temp_buffer[26]), 
         .D(n22432), .Z(MISOb_N_858[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i28_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[27]), .C(temp_buffer[27]), 
         .D(n22432), .Z(MISOb_N_858[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i29_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[28]), .C(temp_buffer[28]), 
         .D(n22432), .Z(MISOb_N_858[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i30_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[29]), .C(temp_buffer[29]), 
         .D(n22432), .Z(MISOb_N_858[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i31_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[30]), .C(temp_buffer[30]), 
         .D(n22432), .Z(MISOb_N_858[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_19 (.A0(recv_buffer[93]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[94]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18821), .COUT(n18822));
    defparam add_15368_19.INIT0 = 16'hf555;
    defparam add_15368_19.INIT1 = 16'hf555;
    defparam add_15368_19.INJECT1_0 = "NO";
    defparam add_15368_19.INJECT1_1 = "NO";
    LUT4 mux_9_i32_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[31]), .C(temp_buffer[31]), 
         .D(n22432), .Z(MISOb_N_858[31])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i32_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_17 (.A0(recv_buffer[91]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[92]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18820), .COUT(n18821));
    defparam add_15368_17.INIT0 = 16'hf555;
    defparam add_15368_17.INIT1 = 16'hf555;
    defparam add_15368_17.INJECT1_0 = "NO";
    defparam add_15368_17.INJECT1_1 = "NO";
    LUT4 mux_9_i33_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[32]), .C(temp_buffer[32]), 
         .D(n22432), .Z(MISOb_N_858[32])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i33_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i34_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[33]), .C(temp_buffer[33]), 
         .D(n22432), .Z(MISOb_N_858[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i35_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[34]), .C(temp_buffer[34]), 
         .D(n22432), .Z(MISOb_N_858[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i36_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[35]), .C(temp_buffer[35]), 
         .D(n22432), .Z(MISOb_N_858[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_15 (.A0(recv_buffer[89]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[90]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18819), .COUT(n18820));
    defparam add_15368_15.INIT0 = 16'hf555;
    defparam add_15368_15.INIT1 = 16'hf555;
    defparam add_15368_15.INJECT1_0 = "NO";
    defparam add_15368_15.INJECT1_1 = "NO";
    CCU2D add_15368_13 (.A0(recv_buffer[87]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[88]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18818), .COUT(n18819));
    defparam add_15368_13.INIT0 = 16'hf555;
    defparam add_15368_13.INIT1 = 16'h0aaa;
    defparam add_15368_13.INJECT1_0 = "NO";
    defparam add_15368_13.INJECT1_1 = "NO";
    LUT4 mux_9_i37_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[36]), .C(temp_buffer[36]), 
         .D(n22432), .Z(MISOb_N_858[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_11 (.A0(recv_buffer[85]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[86]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18817), .COUT(n18818));
    defparam add_15368_11.INIT0 = 16'h0aaa;
    defparam add_15368_11.INIT1 = 16'hf555;
    defparam add_15368_11.INJECT1_0 = "NO";
    defparam add_15368_11.INJECT1_1 = "NO";
    LUT4 mux_9_i38_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[37]), .C(temp_buffer[37]), 
         .D(n22432), .Z(MISOb_N_858[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15382_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18608), 
          .S0(n3496));
    defparam add_15382_cout.INIT0 = 16'h0000;
    defparam add_15382_cout.INIT1 = 16'h0000;
    defparam add_15382_cout.INJECT1_0 = "NO";
    defparam add_15382_cout.INJECT1_1 = "NO";
    CCU2D add_15382_16 (.A0(recv_buffer[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[32]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18607), .COUT(n18608));
    defparam add_15382_16.INIT0 = 16'h5aaa;
    defparam add_15382_16.INIT1 = 16'h0aaa;
    defparam add_15382_16.INJECT1_0 = "NO";
    defparam add_15382_16.INJECT1_1 = "NO";
    CCU2D add_15382_14 (.A0(recv_buffer[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18606), .COUT(n18607));
    defparam add_15382_14.INIT0 = 16'h5aaa;
    defparam add_15382_14.INIT1 = 16'h5aaa;
    defparam add_15382_14.INJECT1_0 = "NO";
    defparam add_15382_14.INJECT1_1 = "NO";
    LUT4 mux_9_i39_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[38]), .C(temp_buffer[38]), 
         .D(n22432), .Z(MISOb_N_858[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i40_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[39]), .C(temp_buffer[39]), 
         .D(n22432), .Z(MISOb_N_858[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i41_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[40]), .C(temp_buffer[40]), 
         .D(n22432), .Z(MISOb_N_858[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i42_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[41]), .C(temp_buffer[41]), 
         .D(n22432), .Z(MISOb_N_858[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15382_12 (.A0(recv_buffer[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18605), .COUT(n18606));
    defparam add_15382_12.INIT0 = 16'h5aaa;
    defparam add_15382_12.INIT1 = 16'h5aaa;
    defparam add_15382_12.INJECT1_0 = "NO";
    defparam add_15382_12.INJECT1_1 = "NO";
    LUT4 mux_9_i43_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[42]), .C(temp_buffer[42]), 
         .D(n22432), .Z(MISOb_N_858[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_9 (.A0(recv_buffer[83]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[84]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18816), .COUT(n18817));
    defparam add_15368_9.INIT0 = 16'h0aaa;
    defparam add_15368_9.INIT1 = 16'h0aaa;
    defparam add_15368_9.INJECT1_0 = "NO";
    defparam add_15368_9.INJECT1_1 = "NO";
    LUT4 mux_9_i44_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[43]), .C(temp_buffer[43]), 
         .D(n22432), .Z(MISOb_N_858[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i45_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[44]), .C(temp_buffer[44]), 
         .D(n22432), .Z(MISOb_N_858[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i46_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[45]), .C(temp_buffer[45]), 
         .D(n22432), .Z(MISOb_N_858[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15382_10 (.A0(recv_buffer[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18604), .COUT(n18605));
    defparam add_15382_10.INIT0 = 16'h5555;
    defparam add_15382_10.INIT1 = 16'h5aaa;
    defparam add_15382_10.INJECT1_0 = "NO";
    defparam add_15382_10.INJECT1_1 = "NO";
    LUT4 mux_9_i47_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[46]), .C(temp_buffer[46]), 
         .D(n22432), .Z(MISOb_N_858[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i48_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[47]), .C(temp_buffer[47]), 
         .D(n22432), .Z(MISOb_N_858[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i49_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[48]), .C(temp_buffer[48]), 
         .D(n22432), .Z(MISOb_N_858[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_7 (.A0(recv_buffer[81]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[82]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18815), .COUT(n18816));
    defparam add_15368_7.INIT0 = 16'hf555;
    defparam add_15368_7.INIT1 = 16'hf555;
    defparam add_15368_7.INJECT1_0 = "NO";
    defparam add_15368_7.INJECT1_1 = "NO";
    CCU2D add_15368_5 (.A0(recv_buffer[79]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[80]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18814), .COUT(n18815));
    defparam add_15368_5.INIT0 = 16'h0aaa;
    defparam add_15368_5.INIT1 = 16'hf555;
    defparam add_15368_5.INJECT1_0 = "NO";
    defparam add_15368_5.INJECT1_1 = "NO";
    CCU2D add_15382_8 (.A0(recv_buffer[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18603), .COUT(n18604));
    defparam add_15382_8.INIT0 = 16'h5aaa;
    defparam add_15382_8.INIT1 = 16'h5aaa;
    defparam add_15382_8.INJECT1_0 = "NO";
    defparam add_15382_8.INJECT1_1 = "NO";
    LUT4 mux_9_i50_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[49]), .C(temp_buffer[49]), 
         .D(n22432), .Z(MISOb_N_858[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15382_6 (.A0(recv_buffer[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18602), .COUT(n18603));
    defparam add_15382_6.INIT0 = 16'h5555;
    defparam add_15382_6.INIT1 = 16'h5555;
    defparam add_15382_6.INJECT1_0 = "NO";
    defparam add_15382_6.INJECT1_1 = "NO";
    CCU2D add_15368_3 (.A0(recv_buffer[77]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[78]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18813), .COUT(n18814));
    defparam add_15368_3.INIT0 = 16'hf555;
    defparam add_15368_3.INIT1 = 16'hf555;
    defparam add_15368_3.INJECT1_0 = "NO";
    defparam add_15368_3.INJECT1_1 = "NO";
    LUT4 mux_9_i51_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[50]), .C(temp_buffer[50]), 
         .D(n22432), .Z(MISOb_N_858[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i52_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[51]), .C(temp_buffer[51]), 
         .D(n22432), .Z(MISOb_N_858[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i53_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[52]), .C(temp_buffer[52]), 
         .D(n22432), .Z(MISOb_N_858[52])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i53_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i54_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[53]), .C(temp_buffer[53]), 
         .D(n22432), .Z(MISOb_N_858[53])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i54_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i55_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[54]), .C(temp_buffer[54]), 
         .D(n22432), .Z(MISOb_N_858[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i56_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[55]), .C(temp_buffer[55]), 
         .D(n22432), .Z(MISOb_N_858[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i57_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[56]), .C(temp_buffer[56]), 
         .D(n22432), .Z(MISOb_N_858[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i58_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[57]), .C(temp_buffer[57]), 
         .D(n22432), .Z(MISOb_N_858[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i59_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[58]), .C(temp_buffer[58]), 
         .D(n22432), .Z(MISOb_N_858[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i60_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[59]), .C(temp_buffer[59]), 
         .D(n22432), .Z(MISOb_N_858[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i61_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[60]), .C(temp_buffer[60]), 
         .D(n22432), .Z(MISOb_N_858[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i62_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[61]), .C(temp_buffer[61]), 
         .D(n22432), .Z(MISOb_N_858[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i63_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[62]), .C(temp_buffer[62]), 
         .D(n22432), .Z(MISOb_N_858[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i64_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[63]), .C(temp_buffer[63]), 
         .D(n22432), .Z(MISOb_N_858[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15382_4 (.A0(recv_buffer[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18601), .COUT(n18602));
    defparam add_15382_4.INIT0 = 16'h5aaa;
    defparam add_15382_4.INIT1 = 16'h5555;
    defparam add_15382_4.INJECT1_0 = "NO";
    defparam add_15382_4.INJECT1_1 = "NO";
    LUT4 mux_9_i65_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[64]), .C(temp_buffer[64]), 
         .D(n22432), .Z(MISOb_N_858[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i66_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[65]), .C(temp_buffer[65]), 
         .D(n22432), .Z(MISOb_N_858[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i67_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[66]), .C(temp_buffer[66]), 
         .D(n22432), .Z(MISOb_N_858[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15368_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[75]), .B1(recv_buffer[76]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18813));
    defparam add_15368_1.INIT0 = 16'hF000;
    defparam add_15368_1.INIT1 = 16'ha666;
    defparam add_15368_1.INJECT1_0 = "NO";
    defparam add_15368_1.INJECT1_1 = "NO";
    LUT4 mux_9_i68_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[67]), .C(temp_buffer[67]), 
         .D(n22432), .Z(MISOb_N_858[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i69_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[68]), .C(temp_buffer[68]), 
         .D(n22432), .Z(MISOb_N_858[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i70_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[69]), .C(temp_buffer[69]), 
         .D(n22432), .Z(MISOb_N_858[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15382_2 (.A0(recv_buffer[17]), .B0(recv_buffer[16]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18601));
    defparam add_15382_2.INIT0 = 16'h7000;
    defparam add_15382_2.INIT1 = 16'h5aaa;
    defparam add_15382_2.INJECT1_0 = "NO";
    defparam add_15382_2.INJECT1_1 = "NO";
    CCU2D add_15383_21 (.A0(recv_buffer[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18600), .S1(n3472));
    defparam add_15383_21.INIT0 = 16'h5555;
    defparam add_15383_21.INIT1 = 16'h0000;
    defparam add_15383_21.INJECT1_0 = "NO";
    defparam add_15383_21.INJECT1_1 = "NO";
    CCU2D add_15383_19 (.A0(recv_buffer[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18599), .COUT(n18600));
    defparam add_15383_19.INIT0 = 16'hf555;
    defparam add_15383_19.INIT1 = 16'hf555;
    defparam add_15383_19.INJECT1_0 = "NO";
    defparam add_15383_19.INJECT1_1 = "NO";
    CCU2D add_15383_17 (.A0(recv_buffer[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18598), .COUT(n18599));
    defparam add_15383_17.INIT0 = 16'hf555;
    defparam add_15383_17.INIT1 = 16'hf555;
    defparam add_15383_17.INJECT1_0 = "NO";
    defparam add_15383_17.INJECT1_1 = "NO";
    LUT4 mux_9_i71_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[70]), .C(temp_buffer[70]), 
         .D(n22432), .Z(MISOb_N_858[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15383_15 (.A0(recv_buffer[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18597), .COUT(n18598));
    defparam add_15383_15.INIT0 = 16'hf555;
    defparam add_15383_15.INIT1 = 16'hf555;
    defparam add_15383_15.INJECT1_0 = "NO";
    defparam add_15383_15.INJECT1_1 = "NO";
    CCU2D add_15383_13 (.A0(recv_buffer[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18596), .COUT(n18597));
    defparam add_15383_13.INIT0 = 16'hf555;
    defparam add_15383_13.INIT1 = 16'h0aaa;
    defparam add_15383_13.INJECT1_0 = "NO";
    defparam add_15383_13.INJECT1_1 = "NO";
    CCU2D add_15383_11 (.A0(recv_buffer[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18595), .COUT(n18596));
    defparam add_15383_11.INIT0 = 16'h0aaa;
    defparam add_15383_11.INIT1 = 16'hf555;
    defparam add_15383_11.INJECT1_0 = "NO";
    defparam add_15383_11.INJECT1_1 = "NO";
    LUT4 mux_9_i72_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[71]), .C(temp_buffer[71]), 
         .D(n22432), .Z(MISOb_N_858[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i73_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[72]), .C(temp_buffer[72]), 
         .D(n22432), .Z(MISOb_N_858[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15383_9 (.A0(recv_buffer[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18594), .COUT(n18595));
    defparam add_15383_9.INIT0 = 16'h0aaa;
    defparam add_15383_9.INIT1 = 16'h0aaa;
    defparam add_15383_9.INJECT1_0 = "NO";
    defparam add_15383_9.INJECT1_1 = "NO";
    CCU2D add_15383_7 (.A0(recv_buffer[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18593), .COUT(n18594));
    defparam add_15383_7.INIT0 = 16'hf555;
    defparam add_15383_7.INIT1 = 16'hf555;
    defparam add_15383_7.INJECT1_0 = "NO";
    defparam add_15383_7.INJECT1_1 = "NO";
    LUT4 mux_9_i74_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[73]), .C(temp_buffer[73]), 
         .D(n22432), .Z(MISOb_N_858[73])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i74_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15383_5 (.A0(recv_buffer[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18592), .COUT(n18593));
    defparam add_15383_5.INIT0 = 16'h0aaa;
    defparam add_15383_5.INIT1 = 16'hf555;
    defparam add_15383_5.INJECT1_0 = "NO";
    defparam add_15383_5.INJECT1_1 = "NO";
    LUT4 mux_9_i75_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[74]), .C(temp_buffer[74]), 
         .D(n22432), .Z(MISOb_N_858[74])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i75_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i76_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[75]), .C(temp_buffer[75]), 
         .D(n22432), .Z(MISOb_N_858[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15383_3 (.A0(recv_buffer[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18591), .COUT(n18592));
    defparam add_15383_3.INIT0 = 16'hf555;
    defparam add_15383_3.INIT1 = 16'hf555;
    defparam add_15383_3.INJECT1_0 = "NO";
    defparam add_15383_3.INJECT1_1 = "NO";
    LUT4 mux_9_i77_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[76]), .C(temp_buffer[76]), 
         .D(n22432), .Z(MISOb_N_858[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15383_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[12]), .B1(recv_buffer[13]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18591));
    defparam add_15383_1.INIT0 = 16'hF000;
    defparam add_15383_1.INIT1 = 16'ha666;
    defparam add_15383_1.INJECT1_0 = "NO";
    defparam add_15383_1.INJECT1_1 = "NO";
    LUT4 mux_9_i78_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[77]), .C(temp_buffer[77]), 
         .D(n22432), .Z(MISOb_N_858[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i79_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[78]), .C(temp_buffer[78]), 
         .D(n22432), .Z(MISOb_N_858[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i80_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[79]), .C(temp_buffer[79]), 
         .D(n22432), .Z(MISOb_N_858[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i81_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[80]), .C(temp_buffer[80]), 
         .D(n22432), .Z(MISOb_N_858[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i82_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[81]), .C(temp_buffer[81]), 
         .D(n22432), .Z(MISOb_N_858[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3IX speed_set_m2_i0_i0 (.D(recv_buffer[54]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i0.GSR = "DISABLED";
    LUT4 mux_9_i83_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[82]), .C(temp_buffer[82]), 
         .D(n22432), .Z(MISOb_N_858[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i84_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[83]), .C(temp_buffer[83]), 
         .D(n22432), .Z(MISOb_N_858[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i85_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[84]), .C(temp_buffer[84]), 
         .D(n22432), .Z(MISOb_N_858[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3IX speed_set_m1_i0_i0 (.D(recv_buffer[75]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i0.GSR = "DISABLED";
    LUT4 mux_9_i86_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[85]), .C(temp_buffer[85]), 
         .D(n22432), .Z(MISOb_N_858[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i87_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[86]), .C(temp_buffer[86]), 
         .D(n22432), .Z(MISOb_N_858[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i88_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[87]), .C(temp_buffer[87]), 
         .D(n22432), .Z(MISOb_N_858[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i89_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[88]), .C(temp_buffer[88]), 
         .D(n22432), .Z(MISOb_N_858[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i90_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[89]), .C(temp_buffer[89]), 
         .D(n22432), .Z(MISOb_N_858[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i91_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[90]), .C(temp_buffer[90]), 
         .D(n22432), .Z(MISOb_N_858[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i92_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[91]), .C(temp_buffer[91]), 
         .D(n22432), .Z(MISOb_N_858[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i93_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[92]), .C(temp_buffer[92]), 
         .D(n22432), .Z(MISOb_N_858[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i94_3_lut_4_lut_4_lut (.A(n22431), .B(send_buffer[93]), .C(temp_buffer[93]), 
         .D(n22432), .Z(MISOb_N_858[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i95_3_lut_4_lut_4_lut (.A(CSlatched), .B(send_buffer[94]), 
         .C(temp_buffer[94]), .D(n22432), .Z(MISOb_N_858[94])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i95_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i2960_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_853), .C(MISOb_N_858[1]), 
         .D(n21690), .Z(MISOb_N_852)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam i2960_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i2_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[1]), 
         .C(MISOb_N_858[2]), .D(n21690), .Z(send_buffer_95__N_442[1])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i2_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i3_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[2]), 
         .C(MISOb_N_858[3]), .D(n21690), .Z(send_buffer_95__N_442[2])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i3_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i4_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[3]), 
         .C(MISOb_N_858[4]), .D(n21690), .Z(send_buffer_95__N_442[3])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i4_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i5_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[4]), 
         .C(MISOb_N_858[5]), .D(n21690), .Z(send_buffer_95__N_442[4])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i5_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i6_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[5]), 
         .C(MISOb_N_858[6]), .D(n21690), .Z(send_buffer_95__N_442[5])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i6_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i7_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[6]), 
         .C(MISOb_N_858[7]), .D(n21690), .Z(send_buffer_95__N_442[6])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i7_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i8_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[7]), 
         .C(MISOb_N_858[8]), .D(n21690), .Z(send_buffer_95__N_442[7])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i8_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i9_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[8]), 
         .C(MISOb_N_858[9]), .D(n21690), .Z(send_buffer_95__N_442[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i10_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[9]), 
         .C(MISOb_N_858[10]), .D(n21690), .Z(send_buffer_95__N_442[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i11_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[10]), 
         .C(MISOb_N_858[11]), .D(n21690), .Z(send_buffer_95__N_442[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i12_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[11]), 
         .C(MISOb_N_858[12]), .D(n21690), .Z(send_buffer_95__N_442[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i13_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[12]), 
         .C(MISOb_N_858[13]), .D(n21690), .Z(send_buffer_95__N_442[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i14_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[13]), 
         .C(MISOb_N_858[14]), .D(n21690), .Z(send_buffer_95__N_442[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i15_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[14]), 
         .C(MISOb_N_858[15]), .D(n21690), .Z(send_buffer_95__N_442[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i16_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[15]), 
         .C(MISOb_N_858[16]), .D(n21690), .Z(send_buffer_95__N_442[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i17_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[16]), 
         .C(MISOb_N_858[17]), .D(n21690), .Z(send_buffer_95__N_442[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i18_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[17]), 
         .C(MISOb_N_858[18]), .D(n21690), .Z(send_buffer_95__N_442[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i19_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[18]), 
         .C(MISOb_N_858[19]), .D(n21690), .Z(send_buffer_95__N_442[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i20_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[19]), 
         .C(MISOb_N_858[20]), .D(n21690), .Z(send_buffer_95__N_442[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i21_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[20]), 
         .C(MISOb_N_858[21]), .D(n21690), .Z(send_buffer_95__N_442[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i22_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[21]), 
         .C(MISOb_N_858[22]), .D(n21690), .Z(send_buffer_95__N_442[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i23_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[22]), 
         .C(MISOb_N_858[23]), .D(n21690), .Z(send_buffer_95__N_442[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i24_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[23]), 
         .C(MISOb_N_858[24]), .D(n21690), .Z(send_buffer_95__N_442[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i25_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[24]), 
         .C(MISOb_N_858[25]), .D(n21690), .Z(send_buffer_95__N_442[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i26_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[25]), 
         .C(MISOb_N_858[26]), .D(n21690), .Z(send_buffer_95__N_442[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i27_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[26]), 
         .C(MISOb_N_858[27]), .D(n21690), .Z(send_buffer_95__N_442[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i28_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[27]), 
         .C(MISOb_N_858[28]), .D(n21690), .Z(send_buffer_95__N_442[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i29_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[28]), 
         .C(MISOb_N_858[29]), .D(n21690), .Z(send_buffer_95__N_442[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i30_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[29]), 
         .C(MISOb_N_858[30]), .D(n21690), .Z(send_buffer_95__N_442[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i31_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[30]), 
         .C(MISOb_N_858[31]), .D(n21690), .Z(send_buffer_95__N_442[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3AX CSlatched_118_rep_422 (.D(CS_c), .SP(clkout_c_enable_272), .CK(clkout_c), 
            .Q(n22431));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_118_rep_422.GSR = "DISABLED";
    LUT4 mux_52_i32_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[31]), 
         .C(MISOb_N_858[32]), .D(n21690), .Z(send_buffer_95__N_442[31])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i32_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i33_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[32]), 
         .C(MISOb_N_858[33]), .D(n21690), .Z(send_buffer_95__N_442[32])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i33_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15367_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18695), 
          .S0(n3352));
    defparam add_15367_cout.INIT0 = 16'h0000;
    defparam add_15367_cout.INIT1 = 16'h0000;
    defparam add_15367_cout.INJECT1_0 = "NO";
    defparam add_15367_cout.INJECT1_1 = "NO";
    LUT4 mux_52_i34_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[33]), 
         .C(MISOb_N_858[34]), .D(n21690), .Z(send_buffer_95__N_442[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15367_16 (.A0(recv_buffer[94]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[95]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18694), .COUT(n18695));
    defparam add_15367_16.INIT0 = 16'h5aaa;
    defparam add_15367_16.INIT1 = 16'h0aaa;
    defparam add_15367_16.INJECT1_0 = "NO";
    defparam add_15367_16.INJECT1_1 = "NO";
    CCU2D add_15367_14 (.A0(recv_buffer[92]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[93]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18693), .COUT(n18694));
    defparam add_15367_14.INIT0 = 16'h5aaa;
    defparam add_15367_14.INIT1 = 16'h5aaa;
    defparam add_15367_14.INJECT1_0 = "NO";
    defparam add_15367_14.INJECT1_1 = "NO";
    LUT4 mux_52_i35_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[34]), 
         .C(MISOb_N_858[35]), .D(n21690), .Z(send_buffer_95__N_442[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i36_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[35]), 
         .C(MISOb_N_858[36]), .D(n21690), .Z(send_buffer_95__N_442[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i37_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[36]), 
         .C(MISOb_N_858[37]), .D(n21690), .Z(send_buffer_95__N_442[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15367_12 (.A0(recv_buffer[90]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[91]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18692), .COUT(n18693));
    defparam add_15367_12.INIT0 = 16'h5aaa;
    defparam add_15367_12.INIT1 = 16'h5aaa;
    defparam add_15367_12.INJECT1_0 = "NO";
    defparam add_15367_12.INJECT1_1 = "NO";
    CCU2D add_15367_10 (.A0(recv_buffer[88]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[89]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18691), .COUT(n18692));
    defparam add_15367_10.INIT0 = 16'h5555;
    defparam add_15367_10.INIT1 = 16'h5aaa;
    defparam add_15367_10.INJECT1_0 = "NO";
    defparam add_15367_10.INJECT1_1 = "NO";
    LUT4 mux_52_i38_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[37]), 
         .C(MISOb_N_858[38]), .D(n21690), .Z(send_buffer_95__N_442[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i39_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[38]), 
         .C(MISOb_N_858[39]), .D(n21690), .Z(send_buffer_95__N_442[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i40_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[39]), 
         .C(MISOb_N_858[40]), .D(n21690), .Z(send_buffer_95__N_442[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i41_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[40]), 
         .C(MISOb_N_858[41]), .D(n21690), .Z(send_buffer_95__N_442[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i42_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[41]), 
         .C(MISOb_N_858[42]), .D(n21690), .Z(send_buffer_95__N_442[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i43_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[42]), 
         .C(MISOb_N_858[43]), .D(n21690), .Z(send_buffer_95__N_442[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i44_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[43]), 
         .C(MISOb_N_858[44]), .D(n21690), .Z(send_buffer_95__N_442[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i45_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[44]), 
         .C(MISOb_N_858[45]), .D(n21690), .Z(send_buffer_95__N_442[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i46_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[45]), 
         .C(MISOb_N_858[46]), .D(n21690), .Z(send_buffer_95__N_442[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i47_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[46]), 
         .C(MISOb_N_858[47]), .D(n21690), .Z(send_buffer_95__N_442[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i48_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[47]), 
         .C(MISOb_N_858[48]), .D(n21690), .Z(send_buffer_95__N_442[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i49_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[48]), 
         .C(MISOb_N_858[49]), .D(n21690), .Z(send_buffer_95__N_442[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i50_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[49]), 
         .C(MISOb_N_858[50]), .D(n21690), .Z(send_buffer_95__N_442[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i51_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[50]), 
         .C(MISOb_N_858[51]), .D(n21690), .Z(send_buffer_95__N_442[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i52_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[51]), 
         .C(MISOb_N_858[52]), .D(n21690), .Z(send_buffer_95__N_442[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i53_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[52]), 
         .C(MISOb_N_858[53]), .D(n21690), .Z(send_buffer_95__N_442[52])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i53_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i54_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[53]), 
         .C(MISOb_N_858[54]), .D(n21690), .Z(send_buffer_95__N_442[53])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i54_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i55_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[54]), 
         .C(MISOb_N_858[55]), .D(n21690), .Z(send_buffer_95__N_442[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i56_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[55]), 
         .C(MISOb_N_858[56]), .D(n21690), .Z(send_buffer_95__N_442[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i57_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[56]), 
         .C(MISOb_N_858[57]), .D(n21690), .Z(send_buffer_95__N_442[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i58_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[57]), 
         .C(MISOb_N_858[58]), .D(n21690), .Z(send_buffer_95__N_442[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i59_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[58]), 
         .C(MISOb_N_858[59]), .D(n21690), .Z(send_buffer_95__N_442[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i60_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[59]), 
         .C(MISOb_N_858[60]), .D(n21690), .Z(send_buffer_95__N_442[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15367_8 (.A0(recv_buffer[86]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[87]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18690), .COUT(n18691));
    defparam add_15367_8.INIT0 = 16'h5aaa;
    defparam add_15367_8.INIT1 = 16'h5aaa;
    defparam add_15367_8.INJECT1_0 = "NO";
    defparam add_15367_8.INJECT1_1 = "NO";
    LUT4 mux_52_i61_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[60]), 
         .C(MISOb_N_858[61]), .D(n21690), .Z(send_buffer_95__N_442[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i62_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[61]), 
         .C(MISOb_N_858[62]), .D(n21690), .Z(send_buffer_95__N_442[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15367_6 (.A0(recv_buffer[84]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[85]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18689), .COUT(n18690));
    defparam add_15367_6.INIT0 = 16'h5555;
    defparam add_15367_6.INIT1 = 16'h5555;
    defparam add_15367_6.INJECT1_0 = "NO";
    defparam add_15367_6.INJECT1_1 = "NO";
    LUT4 mux_52_i63_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[62]), 
         .C(MISOb_N_858[63]), .D(n21690), .Z(send_buffer_95__N_442[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i64_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[63]), 
         .C(MISOb_N_858[64]), .D(n21690), .Z(send_buffer_95__N_442[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15367_4 (.A0(recv_buffer[82]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[83]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18688), .COUT(n18689));
    defparam add_15367_4.INIT0 = 16'h5aaa;
    defparam add_15367_4.INIT1 = 16'h5555;
    defparam add_15367_4.INJECT1_0 = "NO";
    defparam add_15367_4.INJECT1_1 = "NO";
    LUT4 mux_52_i65_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[64]), 
         .C(MISOb_N_858[65]), .D(n21690), .Z(send_buffer_95__N_442[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i66_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[65]), 
         .C(MISOb_N_858[66]), .D(n21690), .Z(send_buffer_95__N_442[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15367_2 (.A0(recv_buffer[80]), .B0(recv_buffer[79]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[81]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18688));
    defparam add_15367_2.INIT0 = 16'h7000;
    defparam add_15367_2.INIT1 = 16'h5aaa;
    defparam add_15367_2.INJECT1_0 = "NO";
    defparam add_15367_2.INJECT1_1 = "NO";
    LUT4 mux_52_i67_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[66]), 
         .C(MISOb_N_858[67]), .D(n21690), .Z(send_buffer_95__N_442[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i68_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[67]), 
         .C(MISOb_N_858[68]), .D(n21690), .Z(send_buffer_95__N_442[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i69_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[68]), 
         .C(MISOb_N_858[69]), .D(n21690), .Z(send_buffer_95__N_442[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i70_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[69]), 
         .C(MISOb_N_858[70]), .D(n21690), .Z(send_buffer_95__N_442[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i71_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[70]), 
         .C(MISOb_N_858[71]), .D(n21690), .Z(send_buffer_95__N_442[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i72_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[71]), 
         .C(MISOb_N_858[72]), .D(n21690), .Z(send_buffer_95__N_442[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i73_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[72]), 
         .C(MISOb_N_858[73]), .D(n21690), .Z(send_buffer_95__N_442[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i74_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[73]), 
         .C(MISOb_N_858[74]), .D(n21690), .Z(send_buffer_95__N_442[73])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i74_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i75_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[74]), 
         .C(MISOb_N_858[75]), .D(n21690), .Z(send_buffer_95__N_442[74])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i75_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i76_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[75]), 
         .C(MISOb_N_858[76]), .D(n21690), .Z(send_buffer_95__N_442[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i77_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[76]), 
         .C(MISOb_N_858[77]), .D(n21690), .Z(send_buffer_95__N_442[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i78_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[77]), 
         .C(MISOb_N_858[78]), .D(n21690), .Z(send_buffer_95__N_442[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i79_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[78]), 
         .C(MISOb_N_858[79]), .D(n21690), .Z(send_buffer_95__N_442[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i80_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[79]), 
         .C(MISOb_N_858[80]), .D(n21690), .Z(send_buffer_95__N_442[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i81_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[80]), 
         .C(MISOb_N_858[81]), .D(n21690), .Z(send_buffer_95__N_442[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i82_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[81]), 
         .C(MISOb_N_858[82]), .D(n21690), .Z(send_buffer_95__N_442[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i83_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[82]), 
         .C(MISOb_N_858[83]), .D(n21690), .Z(send_buffer_95__N_442[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i84_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[83]), 
         .C(MISOb_N_858[84]), .D(n21690), .Z(send_buffer_95__N_442[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i85_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[84]), 
         .C(MISOb_N_858[85]), .D(n21690), .Z(send_buffer_95__N_442[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i86_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[85]), 
         .C(MISOb_N_858[86]), .D(n21690), .Z(send_buffer_95__N_442[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i87_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[86]), 
         .C(MISOb_N_858[87]), .D(n21690), .Z(send_buffer_95__N_442[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i88_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[87]), 
         .C(MISOb_N_858[88]), .D(n21690), .Z(send_buffer_95__N_442[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i89_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[88]), 
         .C(MISOb_N_858[89]), .D(n21690), .Z(send_buffer_95__N_442[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i90_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[89]), 
         .C(MISOb_N_858[90]), .D(n21690), .Z(send_buffer_95__N_442[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i91_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[90]), 
         .C(MISOb_N_858[91]), .D(n21690), .Z(send_buffer_95__N_442[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i92_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[91]), 
         .C(MISOb_N_858[92]), .D(n21690), .Z(send_buffer_95__N_442[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i93_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[92]), 
         .C(MISOb_N_858[93]), .D(n21690), .Z(send_buffer_95__N_442[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i94_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[93]), 
         .C(MISOb_N_858[94]), .D(n21690), .Z(send_buffer_95__N_442[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    FD1P3JX speed_set_m4_i0_i9 (.D(recv_buffer[21]), .SP(clkout_c_enable_350), 
            .PD(n14152), .CK(clkout_c), .Q(speed_set_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i9.GSR = "DISABLED";
    LUT4 mux_52_i95_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[94]), 
         .C(n21662), .D(n21690), .Z(send_buffer_95__N_442[94])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i95_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i143_2_lut_rep_359_3_lut_3_lut (.A(CSlatched), .B(SCKlatched), 
         .C(SCKold), .Z(n21672)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam i143_2_lut_rep_359_3_lut_3_lut.init = 16'h1010;
    FD1P3IX speed_set_m4_i0_i18 (.D(recv_buffer[30]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i18.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i10 (.D(recv_buffer[22]), .SP(clkout_c_enable_350), 
            .PD(n14152), .CK(clkout_c), .Q(speed_set_m4[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i10.GSR = "DISABLED";
    CCU2D add_15384_21 (.A0(recv_buffer[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18794), .S1(n3424));
    defparam add_15384_21.INIT0 = 16'h5555;
    defparam add_15384_21.INIT1 = 16'h0000;
    defparam add_15384_21.INJECT1_0 = "NO";
    defparam add_15384_21.INJECT1_1 = "NO";
    CCU2D add_15384_19 (.A0(recv_buffer[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18793), .COUT(n18794));
    defparam add_15384_19.INIT0 = 16'hf555;
    defparam add_15384_19.INIT1 = 16'hf555;
    defparam add_15384_19.INJECT1_0 = "NO";
    defparam add_15384_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_386 (.A(enable_m4), .B(free_m4), .Z(n21699)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_386.init = 16'h2222;
    LUT4 i17539_3_lut_4_lut (.A(enable_m4), .B(free_m4), .C(hallsense_m4[2]), 
         .D(hallsense_m4[0]), .Z(n19826)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17539_3_lut_4_lut.init = 16'hfddf;
    CCU2D add_15384_17 (.A0(recv_buffer[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18792), .COUT(n18793));
    defparam add_15384_17.INIT0 = 16'hf555;
    defparam add_15384_17.INIT1 = 16'hf555;
    defparam add_15384_17.INJECT1_0 = "NO";
    defparam add_15384_17.INJECT1_1 = "NO";
    CCU2D add_15384_15 (.A0(recv_buffer[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18791), .COUT(n18792));
    defparam add_15384_15.INIT0 = 16'hf555;
    defparam add_15384_15.INIT1 = 16'hf555;
    defparam add_15384_15.INJECT1_0 = "NO";
    defparam add_15384_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_391 (.A(enable_m3), .B(free_m3), .Z(n21704)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_391.init = 16'h2222;
    CCU2D add_15384_13 (.A0(recv_buffer[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18790), .COUT(n18791));
    defparam add_15384_13.INIT0 = 16'hf555;
    defparam add_15384_13.INIT1 = 16'h0aaa;
    defparam add_15384_13.INJECT1_0 = "NO";
    defparam add_15384_13.INJECT1_1 = "NO";
    CCU2D add_15384_11 (.A0(recv_buffer[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18789), .COUT(n18790));
    defparam add_15384_11.INIT0 = 16'h0aaa;
    defparam add_15384_11.INIT1 = 16'hf555;
    defparam add_15384_11.INJECT1_0 = "NO";
    defparam add_15384_11.INJECT1_1 = "NO";
    LUT4 i17528_3_lut_4_lut (.A(enable_m3), .B(free_m3), .C(hallsense_m3[2]), 
         .D(hallsense_m3[0]), .Z(n19845)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17528_3_lut_4_lut.init = 16'hfddf;
    CCU2D add_15384_9 (.A0(recv_buffer[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18788), .COUT(n18789));
    defparam add_15384_9.INIT0 = 16'h0aaa;
    defparam add_15384_9.INIT1 = 16'h0aaa;
    defparam add_15384_9.INJECT1_0 = "NO";
    defparam add_15384_9.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_393 (.A(CSlatched), .B(CSold), .C(n22435), .Z(clkout_c_enable_350)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i2_3_lut_rep_393.init = 16'h8080;
    LUT4 i11643_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22435), .D(enable_m1_N_819), 
         .Z(n14212)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11643_2_lut_4_lut.init = 16'h0080;
    LUT4 i11623_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22435), .D(enable_m2_N_827), 
         .Z(n14192)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11623_2_lut_4_lut.init = 16'h0080;
    FD1P3IX speed_set_m4_i0_i19 (.D(recv_buffer[31]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i19.GSR = "DISABLED";
    LUT4 i11603_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22435), .D(enable_m3_N_834), 
         .Z(n14172)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11603_2_lut_4_lut.init = 16'h0080;
    LUT4 i11583_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22435), .D(enable_m4_N_841), 
         .Z(n14152)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11583_2_lut_4_lut.init = 16'h0080;
    CCU2D add_15384_7 (.A0(recv_buffer[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18787), .COUT(n18788));
    defparam add_15384_7.INIT0 = 16'hf555;
    defparam add_15384_7.INIT1 = 16'hf555;
    defparam add_15384_7.INJECT1_0 = "NO";
    defparam add_15384_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_398 (.A(enable_m2), .B(free_m2), .Z(n21711)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_398.init = 16'h2222;
    LUT4 i17518_3_lut_4_lut (.A(enable_m2), .B(free_m2), .C(hallsense_m2[2]), 
         .D(hallsense_m2[0]), .Z(n19830)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17518_3_lut_4_lut.init = 16'hfddf;
    FD1P3IX speed_set_m1_i0_i1 (.D(recv_buffer[76]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i2 (.D(recv_buffer[77]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i3 (.D(recv_buffer[78]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i4 (.D(recv_buffer[79]), .SP(clkout_c_enable_350), 
            .PD(n14212), .CK(clkout_c), .Q(speed_set_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i5 (.D(recv_buffer[80]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i6 (.D(recv_buffer[81]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i7 (.D(recv_buffer[82]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i8 (.D(recv_buffer[83]), .SP(clkout_c_enable_350), 
            .PD(n14212), .CK(clkout_c), .Q(speed_set_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i9 (.D(recv_buffer[84]), .SP(clkout_c_enable_350), 
            .PD(n14212), .CK(clkout_c), .Q(speed_set_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i10 (.D(recv_buffer[85]), .SP(clkout_c_enable_350), 
            .PD(n14212), .CK(clkout_c), .Q(speed_set_m1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i11 (.D(recv_buffer[86]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i12 (.D(recv_buffer[87]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i13 (.D(recv_buffer[88]), .SP(clkout_c_enable_350), 
            .PD(n14212), .CK(clkout_c), .Q(speed_set_m1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i14 (.D(recv_buffer[89]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i15 (.D(recv_buffer[90]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i16 (.D(recv_buffer[91]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i17 (.D(recv_buffer[92]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i18 (.D(recv_buffer[93]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i19 (.D(recv_buffer[94]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i20 (.D(recv_buffer[95]), .SP(clkout_c_enable_350), 
            .CD(n14212), .CK(clkout_c), .Q(speed_set_m1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i1 (.D(recv_buffer[55]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i2 (.D(recv_buffer[56]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i3 (.D(recv_buffer[57]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i4 (.D(recv_buffer[58]), .SP(clkout_c_enable_350), 
            .PD(n14192), .CK(clkout_c), .Q(speed_set_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i5 (.D(recv_buffer[59]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i6 (.D(recv_buffer[60]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i7 (.D(recv_buffer[61]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i8 (.D(recv_buffer[62]), .SP(clkout_c_enable_350), 
            .PD(n14192), .CK(clkout_c), .Q(speed_set_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i9 (.D(recv_buffer[63]), .SP(clkout_c_enable_350), 
            .PD(n14192), .CK(clkout_c), .Q(speed_set_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i10 (.D(recv_buffer[64]), .SP(clkout_c_enable_350), 
            .PD(n14192), .CK(clkout_c), .Q(speed_set_m2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i11 (.D(recv_buffer[65]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i12 (.D(recv_buffer[66]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i13 (.D(recv_buffer[67]), .SP(clkout_c_enable_350), 
            .PD(n14192), .CK(clkout_c), .Q(speed_set_m2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i14 (.D(recv_buffer[68]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i15 (.D(recv_buffer[69]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i16 (.D(recv_buffer[70]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i17 (.D(recv_buffer[71]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i18 (.D(recv_buffer[72]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i19 (.D(recv_buffer[73]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i19.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_402 (.A(enable_m1), .B(free_m1), .Z(n21715)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_402.init = 16'h2222;
    FD1P3IX speed_set_m2_i0_i20 (.D(recv_buffer[74]), .SP(clkout_c_enable_350), 
            .CD(n14192), .CK(clkout_c), .Q(speed_set_m2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i1 (.D(recv_buffer[34]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i1.GSR = "DISABLED";
    LUT4 i17508_3_lut_4_lut (.A(enable_m1), .B(free_m1), .C(hallsense_m1[2]), 
         .D(hallsense_m1[0]), .Z(n19843)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17508_3_lut_4_lut.init = 16'hfddf;
    FD1P3IX speed_set_m3_i0_i2 (.D(recv_buffer[35]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i3 (.D(recv_buffer[36]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i4 (.D(recv_buffer[37]), .SP(clkout_c_enable_350), 
            .PD(n14172), .CK(clkout_c), .Q(speed_set_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i5 (.D(recv_buffer[38]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i6 (.D(recv_buffer[39]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i7 (.D(recv_buffer[40]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i8 (.D(recv_buffer[41]), .SP(clkout_c_enable_350), 
            .PD(n14172), .CK(clkout_c), .Q(speed_set_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i9 (.D(recv_buffer[42]), .SP(clkout_c_enable_350), 
            .PD(n14172), .CK(clkout_c), .Q(speed_set_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i10 (.D(recv_buffer[43]), .SP(clkout_c_enable_350), 
            .PD(n14172), .CK(clkout_c), .Q(speed_set_m3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i11 (.D(recv_buffer[44]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i12 (.D(recv_buffer[45]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i13 (.D(recv_buffer[46]), .SP(clkout_c_enable_350), 
            .PD(n14172), .CK(clkout_c), .Q(speed_set_m3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i14 (.D(recv_buffer[47]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i15 (.D(recv_buffer[48]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i16 (.D(recv_buffer[49]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i17 (.D(recv_buffer[50]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i18 (.D(recv_buffer[51]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i19 (.D(recv_buffer[52]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i20 (.D(recv_buffer[53]), .SP(clkout_c_enable_350), 
            .CD(n14172), .CK(clkout_c), .Q(speed_set_m3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i1 (.D(recv_buffer[13]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i2 (.D(recv_buffer[14]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i3 (.D(recv_buffer[15]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i4 (.D(recv_buffer[16]), .SP(clkout_c_enable_350), 
            .PD(n14152), .CK(clkout_c), .Q(speed_set_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i4.GSR = "DISABLED";
    FD1P3AX CSold_116_rep_423 (.D(n22431), .SP(clkout_c_enable_341), .CK(clkout_c), 
            .Q(n22432));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_116_rep_423.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i5 (.D(recv_buffer[17]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i5.GSR = "DISABLED";
    LUT4 i13_4_lut_adj_193 (.A(recv_buffer[32]), .B(recv_buffer[31]), .C(recv_buffer[21]), 
         .D(recv_buffer[16]), .Z(n34_adj_2417)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_193.init = 16'hfffe;
    FD1P3IX speed_set_m4_i0_i6 (.D(recv_buffer[18]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i20 (.D(recv_buffer[32]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i11 (.D(recv_buffer[23]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i12 (.D(recv_buffer[24]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i13 (.D(recv_buffer[25]), .SP(clkout_c_enable_350), 
            .PD(n14152), .CK(clkout_c), .Q(speed_set_m4[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i7 (.D(recv_buffer[19]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i7.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i14 (.D(recv_buffer[26]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i15 (.D(recv_buffer[27]), .SP(clkout_c_enable_350), 
            .CD(n14152), .CK(clkout_c), .Q(speed_set_m4[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i15.GSR = "DISABLED";
    CCU2D add_15384_5 (.A0(recv_buffer[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18786), .COUT(n18787));
    defparam add_15384_5.INIT0 = 16'h0aaa;
    defparam add_15384_5.INIT1 = 16'hf555;
    defparam add_15384_5.INJECT1_0 = "NO";
    defparam add_15384_5.INJECT1_1 = "NO";
    CCU2D add_15384_3 (.A0(recv_buffer[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18785), .COUT(n18786));
    defparam add_15384_3.INIT0 = 16'hf555;
    defparam add_15384_3.INIT1 = 16'hf555;
    defparam add_15384_3.INJECT1_0 = "NO";
    defparam add_15384_3.INJECT1_1 = "NO";
    CCU2D add_15384_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[33]), .B1(recv_buffer[34]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18785));
    defparam add_15384_1.INIT0 = 16'hF000;
    defparam add_15384_1.INIT1 = 16'ha666;
    defparam add_15384_1.INJECT1_0 = "NO";
    defparam add_15384_1.INJECT1_1 = "NO";
    PFUMX MISO_I_0 (.BLUT(n5170), .ALUT(MISOb_N_857), .C0(n22435), .Z(MISO_N_862)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;
    
endmodule
//
// Verilog Description of module AVG_SPEED_U9
//

module AVG_SPEED_U9 (\speed_avg_m3[0] , clk_1mhz, \speed_m3[0] , GND_net, 
            \speed_avg_m3[1] , \speed_m3[1] , \speed_avg_m3[2] , \speed_m3[2] , 
            \speed_avg_m3[3] , \speed_m3[3] , \speed_avg_m3[4] , \speed_m3[4] , 
            \speed_avg_m3[5] , \speed_m3[5] , \speed_avg_m3[6] , \speed_m3[6] , 
            \speed_avg_m3[7] , \speed_m3[7] , \speed_avg_m3[8] , \speed_m3[8] , 
            \speed_avg_m3[9] , \speed_m3[9] , \speed_avg_m3[10] , \speed_m3[10] , 
            \speed_avg_m3[11] , \speed_m3[11] , \speed_avg_m3[12] , \speed_m3[12] , 
            \speed_avg_m3[13] , \speed_m3[13] , \speed_avg_m3[14] , \speed_m3[14] , 
            \speed_avg_m3[15] , \speed_m3[15] , \speed_avg_m3[16] , \speed_m3[16] , 
            \speed_avg_m3[17] , \speed_m3[17] , \speed_avg_m3[18] , \speed_m3[18] , 
            \speed_avg_m3[19] , \speed_m3[19] );
    output \speed_avg_m3[0] ;
    input clk_1mhz;
    input \speed_m3[0] ;
    input GND_net;
    output \speed_avg_m3[1] ;
    input \speed_m3[1] ;
    output \speed_avg_m3[2] ;
    input \speed_m3[2] ;
    output \speed_avg_m3[3] ;
    input \speed_m3[3] ;
    output \speed_avg_m3[4] ;
    input \speed_m3[4] ;
    output \speed_avg_m3[5] ;
    input \speed_m3[5] ;
    output \speed_avg_m3[6] ;
    input \speed_m3[6] ;
    output \speed_avg_m3[7] ;
    input \speed_m3[7] ;
    output \speed_avg_m3[8] ;
    input \speed_m3[8] ;
    output \speed_avg_m3[9] ;
    input \speed_m3[9] ;
    output \speed_avg_m3[10] ;
    input \speed_m3[10] ;
    output \speed_avg_m3[11] ;
    input \speed_m3[11] ;
    output \speed_avg_m3[12] ;
    input \speed_m3[12] ;
    output \speed_avg_m3[13] ;
    input \speed_m3[13] ;
    output \speed_avg_m3[14] ;
    input \speed_m3[14] ;
    output \speed_avg_m3[15] ;
    input \speed_m3[15] ;
    output \speed_avg_m3[16] ;
    input \speed_m3[16] ;
    output \speed_avg_m3[17] ;
    input \speed_m3[17] ;
    output \speed_avg_m3[18] ;
    input \speed_m3[18] ;
    output \speed_avg_m3[19] ;
    input \speed_m3[19] ;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_146;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n18546, n18545, n18544, n20154, n6;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m3[0] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2112__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_146), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112__i0.GSR = "DISABLED";
    CCU2D clk_cnt_2112_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18546), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2112_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2112_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2112_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2112_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18545), .COUT(n18546), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2112_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2112_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2112_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2112_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18544), .COUT(n18545), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2112_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2112_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2112_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2112_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18544), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2112_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2112_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2112_add_4_1.INJECT1_1 = "NO";
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m3[1] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m3[2] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m3[3] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m3[4] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m3[5] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m3[6] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m3[7] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m3[8] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m3[9] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m3[10] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m3[11] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m3[12] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m3[13] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m3[14] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m3[15] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m3[16] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m3[17] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m3[18] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m3[19] ), .SP(clk_1mhz_enable_146), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    LUT4 i17550_4_lut (.A(clk_cnt[0]), .B(n20154), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_146)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17550_4_lut.init = 16'h0004;
    LUT4 i16756_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n20154)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16756_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX clk_cnt_2112__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_146), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2112__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_146), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2112__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_146), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2112__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_146), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2112__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_146), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2112__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_146), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2112__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module AVG_SPEED_U10
//

module AVG_SPEED_U10 (GND_net, \speed_avg_m2[0] , clk_1mhz, \speed_m2[0] , 
            \speed_avg_m2[1] , \speed_m2[1] , \speed_avg_m2[2] , \speed_m2[2] , 
            \speed_avg_m2[3] , \speed_m2[3] , \speed_avg_m2[4] , \speed_m2[4] , 
            \speed_avg_m2[5] , \speed_m2[5] , \speed_avg_m2[6] , \speed_m2[6] , 
            \speed_avg_m2[7] , \speed_m2[7] , \speed_avg_m2[8] , \speed_m2[8] , 
            \speed_avg_m2[9] , \speed_m2[9] , \speed_avg_m2[10] , \speed_m2[10] , 
            \speed_avg_m2[11] , \speed_m2[11] , \speed_avg_m2[12] , \speed_m2[12] , 
            \speed_avg_m2[13] , \speed_m2[13] , \speed_avg_m2[14] , \speed_m2[14] , 
            \speed_avg_m2[15] , \speed_m2[15] , \speed_avg_m2[16] , \speed_m2[16] , 
            \speed_avg_m2[17] , \speed_m2[17] , \speed_avg_m2[18] , \speed_m2[18] , 
            \speed_avg_m2[19] , \speed_m2[19] );
    input GND_net;
    output \speed_avg_m2[0] ;
    input clk_1mhz;
    input \speed_m2[0] ;
    output \speed_avg_m2[1] ;
    input \speed_m2[1] ;
    output \speed_avg_m2[2] ;
    input \speed_m2[2] ;
    output \speed_avg_m2[3] ;
    input \speed_m2[3] ;
    output \speed_avg_m2[4] ;
    input \speed_m2[4] ;
    output \speed_avg_m2[5] ;
    input \speed_m2[5] ;
    output \speed_avg_m2[6] ;
    input \speed_m2[6] ;
    output \speed_avg_m2[7] ;
    input \speed_m2[7] ;
    output \speed_avg_m2[8] ;
    input \speed_m2[8] ;
    output \speed_avg_m2[9] ;
    input \speed_m2[9] ;
    output \speed_avg_m2[10] ;
    input \speed_m2[10] ;
    output \speed_avg_m2[11] ;
    input \speed_m2[11] ;
    output \speed_avg_m2[12] ;
    input \speed_m2[12] ;
    output \speed_avg_m2[13] ;
    input \speed_m2[13] ;
    output \speed_avg_m2[14] ;
    input \speed_m2[14] ;
    output \speed_avg_m2[15] ;
    input \speed_m2[15] ;
    output \speed_avg_m2[16] ;
    input \speed_m2[16] ;
    output \speed_avg_m2[17] ;
    input \speed_m2[17] ;
    output \speed_avg_m2[18] ;
    input \speed_m2[18] ;
    output \speed_avg_m2[19] ;
    input \speed_m2[19] ;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire n18550;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n18549, clk_1mhz_enable_127, n18548, n20132, n6;
    
    CCU2D clk_cnt_2110_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18550), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2110_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2110_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2110_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2110_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18549), .COUT(n18550), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2110_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2110_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2110_add_4_5.INJECT1_1 = "NO";
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m2[0] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    CCU2D clk_cnt_2110_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18548), .COUT(n18549), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2110_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2110_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2110_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2110_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18548), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2110_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2110_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2110_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2110__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_127), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110__i0.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m2[1] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m2[2] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m2[3] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m2[4] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m2[5] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m2[6] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m2[7] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m2[8] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m2[9] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m2[10] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m2[11] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m2[12] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m2[13] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m2[14] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m2[15] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m2[16] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m2[17] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m2[18] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m2[19] ), .SP(clk_1mhz_enable_127), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    LUT4 i17556_4_lut (.A(clk_cnt[4]), .B(n20132), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_127)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17556_4_lut.init = 16'h0004;
    LUT4 i16734_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n20132)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16734_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX clk_cnt_2110__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_127), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2110__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_127), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2110__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_127), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2110__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_127), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2110__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_127), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2110__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_127), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2110__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module AVG_SPEED_U11
//

module AVG_SPEED_U11 (GND_net, \speed_avg_m1[0] , clk_1mhz, \speed_m1[0] , 
            \speed_avg_m1[1] , \speed_m1[1] , \speed_avg_m1[2] , \speed_m1[2] , 
            \speed_avg_m1[3] , \speed_m1[3] , \speed_avg_m1[4] , \speed_m1[4] , 
            \speed_avg_m1[5] , \speed_m1[5] , \speed_avg_m1[6] , \speed_m1[6] , 
            \speed_avg_m1[7] , \speed_m1[7] , \speed_avg_m1[8] , \speed_m1[8] , 
            \speed_avg_m1[9] , \speed_m1[9] , \speed_avg_m1[10] , \speed_m1[10] , 
            \speed_avg_m1[11] , \speed_m1[11] , \speed_avg_m1[12] , \speed_m1[12] , 
            \speed_avg_m1[13] , \speed_m1[13] , \speed_avg_m1[14] , \speed_m1[14] , 
            \speed_avg_m1[15] , \speed_m1[15] , \speed_avg_m1[16] , \speed_m1[16] , 
            \speed_avg_m1[17] , \speed_m1[17] , \speed_avg_m1[18] , \speed_m1[18] , 
            \speed_avg_m1[19] , \speed_m1[19] );
    input GND_net;
    output \speed_avg_m1[0] ;
    input clk_1mhz;
    input \speed_m1[0] ;
    output \speed_avg_m1[1] ;
    input \speed_m1[1] ;
    output \speed_avg_m1[2] ;
    input \speed_m1[2] ;
    output \speed_avg_m1[3] ;
    input \speed_m1[3] ;
    output \speed_avg_m1[4] ;
    input \speed_m1[4] ;
    output \speed_avg_m1[5] ;
    input \speed_m1[5] ;
    output \speed_avg_m1[6] ;
    input \speed_m1[6] ;
    output \speed_avg_m1[7] ;
    input \speed_m1[7] ;
    output \speed_avg_m1[8] ;
    input \speed_m1[8] ;
    output \speed_avg_m1[9] ;
    input \speed_m1[9] ;
    output \speed_avg_m1[10] ;
    input \speed_m1[10] ;
    output \speed_avg_m1[11] ;
    input \speed_m1[11] ;
    output \speed_avg_m1[12] ;
    input \speed_m1[12] ;
    output \speed_avg_m1[13] ;
    input \speed_m1[13] ;
    output \speed_avg_m1[14] ;
    input \speed_m1[14] ;
    output \speed_avg_m1[15] ;
    input \speed_m1[15] ;
    output \speed_avg_m1[16] ;
    input \speed_m1[16] ;
    output \speed_avg_m1[17] ;
    input \speed_m1[17] ;
    output \speed_avg_m1[18] ;
    input \speed_m1[18] ;
    output \speed_avg_m1[19] ;
    input \speed_m1[19] ;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire n18553;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n18554, n18552, clk_1mhz_enable_108, n20130, n6;
    
    CCU2D clk_cnt_2108_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18553), .COUT(n18554), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2108_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2108_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2108_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2108_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18552), .COUT(n18553), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2108_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2108_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2108_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2108_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18552), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2108_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2108_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2108_add_4_1.INJECT1_1 = "NO";
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m1[0] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2108__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_108), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108__i0.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m1[1] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m1[2] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m1[3] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m1[4] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m1[5] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m1[6] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m1[7] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m1[8] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m1[9] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m1[10] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m1[11] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m1[12] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m1[13] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m1[14] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m1[15] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m1[16] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m1[17] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m1[18] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m1[19] ), .SP(clk_1mhz_enable_108), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    LUT4 i17553_4_lut (.A(clk_cnt[0]), .B(n20130), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_108)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17553_4_lut.init = 16'h0004;
    LUT4 i16732_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n20130)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16732_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX clk_cnt_2108__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_108), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2108__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_108), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2108__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_108), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2108__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_108), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2108__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_108), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2108__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_108), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108__i6.GSR = "DISABLED";
    CCU2D clk_cnt_2108_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18554), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2108_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2108_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2108_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2108_add_4_7.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module HALL_U3
//

module HALL_U3 (clk_1mhz, n22430, \speed_m3[0] , hallsense_m3, clkout_c_enable_341, 
            H_A_m3_c, H_B_m3_c, H_C_m3_c, \speed_m3[1] , \speed_m3[2] , 
            \speed_m3[3] , \speed_m3[4] , \speed_m3[5] , \speed_m3[6] , 
            \speed_m3[7] , \speed_m3[8] , \speed_m3[9] , \speed_m3[10] , 
            \speed_m3[11] , \speed_m3[12] , \speed_m3[13] , \speed_m3[14] , 
            \speed_m3[15] , \speed_m3[16] , \speed_m3[17] , \speed_m3[18] , 
            \speed_m3[19] , GND_net);
    input clk_1mhz;
    input n22430;
    output \speed_m3[0] ;
    output [2:0]hallsense_m3;
    input clkout_c_enable_341;
    input H_A_m3_c;
    input H_B_m3_c;
    input H_C_m3_c;
    output \speed_m3[1] ;
    output \speed_m3[2] ;
    output \speed_m3[3] ;
    output \speed_m3[4] ;
    output \speed_m3[5] ;
    output \speed_m3[6] ;
    output \speed_m3[7] ;
    output \speed_m3[8] ;
    output \speed_m3[9] ;
    output \speed_m3[10] ;
    output \speed_m3[11] ;
    output \speed_m3[12] ;
    output \speed_m3[13] ;
    output \speed_m3[14] ;
    output \speed_m3[15] ;
    output \speed_m3[16] ;
    output \speed_m3[17] ;
    output \speed_m3[18] ;
    output \speed_m3[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire stable_counting, clk_1mhz_enable_3, n14384;
    wire [19:0]speedt_19__N_2047;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4597;
    wire [19:0]count_19__N_2067;
    
    wire hall3_lat;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_184, hall3_old, hall1_lat, hall2_lat, hall1_old, 
        hall2_old;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21689;
    wire [6:0]n63;
    
    wire n4, n21670, n19931, n19847, n20120, n20168, n20112, n11461, 
        n20108, n19978, n19806, n11449, stable_counting_N_2129, n21669, 
        n21655, n18476, n18477, n18475, n18474, n18473, n19079, 
        n20026, n19, n24, n20, n21641, n4_adj_2393, n22, n16, 
        n12, n18482, n18481, n18480, n18479, n18478;
    
    FD1P3IX stable_counting_62 (.D(n22430), .SP(clk_1mhz_enable_3), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_2047[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_19__N_2067[0]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2067[0]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m3_c), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m3_c), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m3_c), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 i2508_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21689), .C(stable_count[4]), 
         .D(stable_count[3]), .Z(n63[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2508_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2_3_lut_rep_357 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(n21670)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_357.init = 16'hdede;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .D(n63[1]), 
         .Z(n19931)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 i2485_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2485_1_lut.init = 16'h5555;
    FD1P3AX speed__i2 (.D(speedt_19__N_2047[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2047[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2047[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2047[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2047[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2047[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2047[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2047[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2047[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2047[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2047[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2047[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2047[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2047[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2047[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2047[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2047[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2047[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2047[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(count_19__N_2067[1]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2067[2]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2067[3]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2067[4]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2067[5]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2067[6]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2067[7]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2067[8]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2067[9]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2067[10]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2067[11]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2067[12]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2067[13]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2067[14]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2067[15]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2067[16]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2067[17]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2067[18]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2067[19]), .CK(clk_1mhz), .CD(n4597), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n19847), .B(n20120), .C(n20168), .D(n20112), .Z(n11461)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0002;
    LUT4 i16722_2_lut (.A(count[11]), .B(count[14]), .Z(n20120)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16722_2_lut.init = 16'heeee;
    LUT4 i16770_4_lut (.A(count[18]), .B(n20108), .C(n19978), .D(count[16]), 
         .Z(n20168)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16770_4_lut.init = 16'hfffe;
    LUT4 i16714_3_lut (.A(count[12]), .B(count[4]), .C(count[15]), .Z(n20112)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16714_3_lut.init = 16'hfefe;
    LUT4 i16710_4_lut (.A(count[5]), .B(count[7]), .C(count[6]), .D(count[17]), 
         .Z(n20108)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16710_4_lut.init = 16'hfffe;
    LUT4 i16581_2_lut (.A(count[1]), .B(count[19]), .Z(n19978)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16581_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(n63[4]), .B(stable_count[0]), .C(n19806), .D(n19931), 
         .Z(n11449)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i2273_2_lut (.A(stable_counting), .B(stable_counting_N_2129), .Z(n4597)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2273_2_lut.init = 16'h8888;
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2067[1]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2067[2]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2067[3]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2067[4]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2067[5]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2067[6]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2067[7]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2067[8]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2067[9]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2067[10]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2067[11]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2067[12]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2067[13]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2067[14]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2067[15]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2067[16]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2067[17]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2067[18]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2067[19]), .SP(clk_1mhz_enable_184), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2047[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2047[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2047[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2047[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2047[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2047[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2047[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2047[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2047[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2047[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2047[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2047[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2047[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2047[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2047[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2047[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2047[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2047[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2047[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11461), .B(n11449), .C(count_19__N_2067[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2047[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i11514_4_lut (.A(n11461), .B(n11449), .C(stable_counting), .D(stable_counting_N_2129), 
         .Z(clk_1mhz_enable_184)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11514_4_lut.init = 16'hcaea;
    LUT4 i2489_2_lut_rep_376 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21689)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2489_2_lut_rep_376.init = 16'h8888;
    LUT4 i2494_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2494_2_lut_3_lut.init = 16'h7878;
    LUT4 i2496_2_lut_rep_356_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21669)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2496_2_lut_rep_356_3_lut.init = 16'h8080;
    LUT4 i2503_2_lut_rep_342_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21655)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2503_2_lut_rep_342_3_lut_4_lut.init = 16'h8000;
    LUT4 i2501_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2501_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18476), 
          .COUT(n18477), .S0(count_19__N_2067[7]), .S1(count_19__N_2067[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18475), 
          .COUT(n18476), .S0(count_19__N_2067[5]), .S1(count_19__N_2067[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18474), 
          .COUT(n18475), .S0(count_19__N_2067[3]), .S1(count_19__N_2067[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18473), 
          .COUT(n18474), .S0(count_19__N_2067[1]), .S1(count_19__N_2067[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18473), 
          .S1(count_19__N_2067[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i17458_4_lut (.A(n19079), .B(n20026), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_3)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17458_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_156 (.A(n19), .B(n19847), .C(n24), .D(n20), .Z(n19079)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_156.init = 16'hfffb;
    LUT4 i1_2_lut_4_lut_adj_157 (.A(n63[6]), .B(n63[3]), .C(n21641), .D(stable_count[0]), 
         .Z(n4_adj_2393)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_2_lut_4_lut_adj_157.init = 16'hfeff;
    LUT4 i16629_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n20026)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16629_4_lut.init = 16'h7bde;
    LUT4 i1_2_lut_4_lut_adj_158 (.A(n63[6]), .B(n63[3]), .C(n21641), .D(n63[2]), 
         .Z(n19806)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_2_lut_4_lut_adj_158.init = 16'hfffe;
    LUT4 i6_2_lut (.A(count[17]), .B(count[11]), .Z(n19)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i11_4_lut (.A(count[5]), .B(n22), .C(n16), .D(count[16]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut (.A(count[14]), .B(count[19]), .C(count[6]), .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i9_4_lut (.A(count[18]), .B(count[12]), .C(count[4]), .D(count[7]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[15]), .B(count[1]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i16748_3_lut (.A(n21670), .B(stable_counting), .C(stable_counting_N_2129), 
         .Z(n14384)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16748_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_159 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_159.init = 16'h7bde;
    LUT4 i2522_3_lut_4_lut (.A(stable_count[4]), .B(n21655), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2522_3_lut_4_lut.init = 16'h7f80;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21641), .SP(stable_counting), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n63[4]), .SP(stable_counting), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(n19931), .B(n63[2]), .C(n63[4]), .D(n4_adj_2393), 
         .Z(stable_counting_N_2129)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i2_4_lut.init = 16'h0002;
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14384), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    LUT4 i2487_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2487_2_lut.init = 16'h6666;
    LUT4 i6_4_lut (.A(count[10]), .B(n12), .C(count[9]), .D(count[2]), 
         .Z(n19847)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[3]), .B(count[8]), .C(count[13]), .D(count[0]), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i2515_2_lut_rep_328_3_lut_4_lut (.A(stable_count[3]), .B(n21669), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21641)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2515_2_lut_rep_328_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18482), 
          .S0(count_19__N_2067[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18481), .COUT(n18482), .S0(count_19__N_2067[17]), .S1(count_19__N_2067[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18480), .COUT(n18481), .S0(count_19__N_2067[15]), .S1(count_19__N_2067[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18479), .COUT(n18480), .S0(count_19__N_2067[13]), .S1(count_19__N_2067[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18478), .COUT(n18479), .S0(count_19__N_2067[11]), .S1(count_19__N_2067[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18477), .COUT(n18478), .S0(count_19__N_2067[9]), .S1(count_19__N_2067[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U1
//

module PWMGENERATOR_U1 (PWM_m2, pwm_clk, free_m2, clkout_c_enable_341, 
            PWMdut_m2, GND_net, hallsense_m2, n21710, enable_m2, n3028, 
            n21712, n2992);
    output PWM_m2;
    input pwm_clk;
    output free_m2;
    input clkout_c_enable_341;
    input [9:0]PWMdut_m2;
    input GND_net;
    input [2:0]hallsense_m2;
    output n21710;
    input enable_m2;
    output n3028;
    output n21712;
    output n2992;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_2176, free_N_2188, n3870, n10, n7, n10_adj_2391, 
        n11438, n9, n17;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    
    wire n16, n14149, n14, n10_adj_2392, n18522, n18521, n18520, 
        n18519, n18518, n18570;
    wire [9:0]n45;
    
    wire n18569, n18568, n18567, n18566;
    
    FD1S3AX PWM_20 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m2)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_2188), .SP(clkout_c_enable_341), .CK(pwm_clk), 
            .Q(free_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i1806_1_lut (.A(n3870), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1806_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(PWMdut_m2[5]), .B(PWMdut_m2[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_2391), .B(PWMdut_m2[9]), .C(PWMdut_m2[8]), 
         .D(PWMdut_m2[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2306_3_lut (.A(n11438), .B(PWMdut_m2[4]), .C(PWMdut_m2[3]), 
         .Z(n10_adj_2391)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2306_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i17491_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n14149)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17491_4_lut.init = 16'h0400;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i6_4_lut (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut.init = 16'hffef;
    LUT4 i17469_4_lut (.A(PWMdut_m2[5]), .B(n14), .C(n10_adj_2392), .D(PWMdut_m2[8]), 
         .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17469_4_lut.init = 16'h0001;
    LUT4 i6_4_lut_adj_154 (.A(PWMdut_m2[9]), .B(PWMdut_m2[3]), .C(PWMdut_m2[4]), 
         .D(n11438), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut_adj_154.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[7]), .Z(n10_adj_2392)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_155 (.A(PWMdut_m2[2]), .B(PWMdut_m2[1]), .C(PWMdut_m2[0]), 
         .Z(n11438)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_155.init = 16'hfefe;
    CCU2D sub_1804_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m2[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18522), .S1(n3870));
    defparam sub_1804_add_2_11.INIT0 = 16'h5999;
    defparam sub_1804_add_2_11.INIT1 = 16'h0000;
    defparam sub_1804_add_2_11.INJECT1_0 = "NO";
    defparam sub_1804_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_9 (.A0(PWMdut_m2[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m2[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18521), 
          .COUT(n18522));
    defparam sub_1804_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1804_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1804_add_2_9.INJECT1_0 = "NO";
    defparam sub_1804_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_7 (.A0(PWMdut_m2[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m2[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18520), 
          .COUT(n18521));
    defparam sub_1804_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1804_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1804_add_2_7.INJECT1_0 = "NO";
    defparam sub_1804_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_5 (.A0(PWMdut_m2[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m2[4]), .C1(n9), .D1(n10), .CIN(n18519), 
          .COUT(n18520));
    defparam sub_1804_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1804_add_2_5.INIT1 = 16'h5999;
    defparam sub_1804_add_2_5.INJECT1_0 = "NO";
    defparam sub_1804_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m2[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m2[2]), .C1(n9), .D1(n10), .CIN(n18518), 
          .COUT(n18519));
    defparam sub_1804_add_2_3.INIT0 = 16'h5999;
    defparam sub_1804_add_2_3.INIT1 = 16'h5999;
    defparam sub_1804_add_2_3.INJECT1_0 = "NO";
    defparam sub_1804_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m2[0]), .C1(n9), .D1(n10), 
          .COUT(n18518));
    defparam sub_1804_add_2_1.INIT0 = 16'h0000;
    defparam sub_1804_add_2_1.INIT1 = 16'h5999;
    defparam sub_1804_add_2_1.INJECT1_0 = "NO";
    defparam sub_1804_add_2_1.INJECT1_1 = "NO";
    CCU2D cnt_2104_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18570), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2104_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2104_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2104_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2104_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18569), 
          .COUT(n18570), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2104_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2104_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2104_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2104_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18568), 
          .COUT(n18569), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2104_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2104_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2104_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2104_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18567), 
          .COUT(n18568), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2104_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2104_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2104_add_4_5.INJECT1_1 = "NO";
    LUT4 i1542_3_lut_rep_397 (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .Z(n21710)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1542_3_lut_rep_397.init = 16'h1414;
    LUT4 i17514_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .D(enable_m2), .Z(n3028)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17514_2_lut_4_lut.init = 16'hebff;
    LUT4 i1512_3_lut_rep_399 (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .Z(n21712)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1512_3_lut_rep_399.init = 16'h1414;
    LUT4 i17511_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .D(enable_m2), .Z(n2992)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17511_2_lut_4_lut.init = 16'hebff;
    CCU2D cnt_2104_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18566), 
          .COUT(n18567), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2104_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2104_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2104_add_4_3.INJECT1_1 = "NO";
    FD1S3IX cnt_2104__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14149), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i0.GSR = "ENABLED";
    CCU2D cnt_2104_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18566), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2104_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2104_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2104_add_4_1.INJECT1_1 = "NO";
    FD1S3IX cnt_2104__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14149), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i1.GSR = "ENABLED";
    FD1S3IX cnt_2104__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14149), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i2.GSR = "ENABLED";
    FD1S3IX cnt_2104__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14149), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i3.GSR = "ENABLED";
    FD1S3IX cnt_2104__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14149), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i4.GSR = "ENABLED";
    FD1S3IX cnt_2104__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14149), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i5.GSR = "ENABLED";
    FD1S3IX cnt_2104__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14149), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i6.GSR = "ENABLED";
    FD1S3IX cnt_2104__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14149), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i7.GSR = "ENABLED";
    FD1S3IX cnt_2104__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14149), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i8.GSR = "ENABLED";
    FD1S3IX cnt_2104__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14149), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2104__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION
//

module COMMUTATION (MB_m4_c_0, clkout_c, MC_m4_c_0, MA_m4_c_0, LED4_c, 
            enable_m4, n3196, n21700, PWM_m4, n3232, n21696, n19826, 
            n21695, free_m4, MA_m4_c_1, n3290, MC_m4_c_1, n3244, 
            MB_m4_c_1, n3208);
    output MB_m4_c_0;
    input clkout_c;
    output MC_m4_c_0;
    output MA_m4_c_0;
    output LED4_c;
    input enable_m4;
    input n3196;
    input n21700;
    input PWM_m4;
    input n3232;
    input n21696;
    input n19826;
    input n21695;
    input free_m4;
    output MA_m4_c_1;
    input n3290;
    output MC_m4_c_1;
    input n3244;
    output MB_m4_c_1;
    input n3208;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_2151, n18968, n18967, n19827, n14105;
    
    FD1S3IX MospairB_i1 (.D(n18968), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MB_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18967), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MC_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19827), .CK(clkout_c), .CD(led1_N_2151), 
            .Q(MA_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14105), .CK(clkout_c), .PD(led1_N_2151), .Q(LED4_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10635_1_lut (.A(enable_m4), .Z(led1_N_2151)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10635_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3196), .B(n21700), .C(PWM_m4), .Z(n18968)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_153 (.A(n3232), .B(n21696), .C(PWM_m4), .Z(n18967)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_153.init = 16'hbfbf;
    LUT4 i17574_3_lut (.A(n19826), .B(PWM_m4), .C(n21695), .Z(n19827)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17574_3_lut.init = 16'hbfbf;
    LUT4 i11518_2_lut (.A(free_m4), .B(LED4_c), .Z(n14105)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11518_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n3290), .CK(clkout_c), .CD(n19826), .Q(MA_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3232), .CK(clkout_c), .CD(n3244), .Q(MC_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3196), .CK(clkout_c), .CD(n3208), .Q(MB_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U2
//

module PWMGENERATOR_U2 (PWM_m1, pwm_clk, free_m1, clkout_c_enable_341, 
            PWMdut_m1, GND_net, hallsense_m1, n21714, enable_m1, n2920, 
            n21716, n2884);
    output PWM_m1;
    input pwm_clk;
    output free_m1;
    input clkout_c_enable_341;
    input [9:0]PWMdut_m1;
    input GND_net;
    input [2:0]hallsense_m1;
    output n21714;
    input enable_m1;
    output n2920;
    output n21716;
    output n2884;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_2176, free_N_2188, n3857, n10, n7, n10_adj_2389, 
        n11436, n9, n17;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    
    wire n16, n14150, n18527, n18526, n18525, n18524, n18523, 
        n14, n10_adj_2390, n18575;
    wire [9:0]n45;
    
    wire n18574, n18573, n18572, n18571;
    
    FD1S3AX PWM_20 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_2188), .SP(clkout_c_enable_341), .CK(pwm_clk), 
            .Q(free_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i1804_1_lut (.A(n3857), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1804_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(PWMdut_m1[5]), .B(PWMdut_m1[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_2389), .B(PWMdut_m1[9]), .C(PWMdut_m1[8]), 
         .D(PWMdut_m1[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2337_3_lut (.A(n11436), .B(PWMdut_m1[4]), .C(PWMdut_m1[3]), 
         .Z(n10_adj_2389)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2337_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i17494_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n14150)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17494_4_lut.init = 16'h0400;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i6_4_lut (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut.init = 16'hffef;
    CCU2D sub_1802_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m1[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18527), .S1(n3857));
    defparam sub_1802_add_2_11.INIT0 = 16'h5999;
    defparam sub_1802_add_2_11.INIT1 = 16'h0000;
    defparam sub_1802_add_2_11.INJECT1_0 = "NO";
    defparam sub_1802_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_9 (.A0(PWMdut_m1[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m1[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18526), 
          .COUT(n18527));
    defparam sub_1802_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1802_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1802_add_2_9.INJECT1_0 = "NO";
    defparam sub_1802_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_7 (.A0(PWMdut_m1[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m1[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18525), 
          .COUT(n18526));
    defparam sub_1802_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1802_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1802_add_2_7.INJECT1_0 = "NO";
    defparam sub_1802_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_5 (.A0(PWMdut_m1[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m1[4]), .C1(n9), .D1(n10), .CIN(n18524), 
          .COUT(n18525));
    defparam sub_1802_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1802_add_2_5.INIT1 = 16'h5999;
    defparam sub_1802_add_2_5.INJECT1_0 = "NO";
    defparam sub_1802_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m1[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m1[2]), .C1(n9), .D1(n10), .CIN(n18523), 
          .COUT(n18524));
    defparam sub_1802_add_2_3.INIT0 = 16'h5999;
    defparam sub_1802_add_2_3.INIT1 = 16'h5999;
    defparam sub_1802_add_2_3.INJECT1_0 = "NO";
    defparam sub_1802_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m1[0]), .C1(n9), .D1(n10), 
          .COUT(n18523));
    defparam sub_1802_add_2_1.INIT0 = 16'h0000;
    defparam sub_1802_add_2_1.INIT1 = 16'h5999;
    defparam sub_1802_add_2_1.INJECT1_0 = "NO";
    defparam sub_1802_add_2_1.INJECT1_1 = "NO";
    LUT4 i17472_4_lut (.A(PWMdut_m1[5]), .B(n14), .C(n10_adj_2390), .D(PWMdut_m1[8]), 
         .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17472_4_lut.init = 16'h0001;
    LUT4 i6_4_lut_adj_151 (.A(PWMdut_m1[9]), .B(PWMdut_m1[3]), .C(PWMdut_m1[4]), 
         .D(n11436), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut_adj_151.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[7]), .Z(n10_adj_2390)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_152 (.A(PWMdut_m1[2]), .B(PWMdut_m1[1]), .C(PWMdut_m1[0]), 
         .Z(n11436)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_152.init = 16'hfefe;
    CCU2D cnt_2103_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18575), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2103_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2103_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2103_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2103_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18574), 
          .COUT(n18575), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2103_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2103_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2103_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2103_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18573), 
          .COUT(n18574), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2103_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2103_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2103_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2103_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18572), 
          .COUT(n18573), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2103_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2103_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2103_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2103_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18571), 
          .COUT(n18572), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2103_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2103_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2103_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2103_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18571), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2103_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2103_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2103_add_4_1.INJECT1_1 = "NO";
    LUT4 i1452_3_lut_rep_401 (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .Z(n21714)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1452_3_lut_rep_401.init = 16'h1414;
    LUT4 i17504_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .D(enable_m1), .Z(n2920)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17504_2_lut_4_lut.init = 16'hebff;
    LUT4 i1422_3_lut_rep_403 (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .Z(n21716)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1422_3_lut_rep_403.init = 16'h1414;
    LUT4 i17501_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .D(enable_m1), .Z(n2884)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17501_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2103__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14150), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i0.GSR = "ENABLED";
    FD1S3IX cnt_2103__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14150), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i1.GSR = "ENABLED";
    FD1S3IX cnt_2103__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14150), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i2.GSR = "ENABLED";
    FD1S3IX cnt_2103__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14150), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i3.GSR = "ENABLED";
    FD1S3IX cnt_2103__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14150), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i4.GSR = "ENABLED";
    FD1S3IX cnt_2103__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14150), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i5.GSR = "ENABLED";
    FD1S3IX cnt_2103__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14150), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i6.GSR = "ENABLED";
    FD1S3IX cnt_2103__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14150), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i7.GSR = "ENABLED";
    FD1S3IX cnt_2103__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14150), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i8.GSR = "ENABLED";
    FD1S3IX cnt_2103__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14150), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2103__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U0
//

module PWMGENERATOR_U0 (PWM_m3, pwm_clk, free_m3, clkout_c_enable_341, 
            PWMdut_m3, GND_net, hallsense_m3, n21703, enable_m3, n3136, 
            n21705, n3100);
    output PWM_m3;
    input pwm_clk;
    output free_m3;
    input clkout_c_enable_341;
    input [9:0]PWMdut_m3;
    input GND_net;
    input [2:0]hallsense_m3;
    output n21703;
    input enable_m3;
    output n3136;
    output n21705;
    output n3100;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_2176, free_N_2188, n3883, n10, n7;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    
    wire n20176, n6, n14148, n20134, n10_adj_2387, n11440, n9, 
        n14, n10_adj_2388, n18517, n18516, n18515, n18514, n18513;
    wire [9:0]n45;
    
    wire n18565, n18564, n18563, n18562, n18561;
    
    FD1S3AX PWM_20 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m3)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_2188), .SP(clkout_c_enable_341), .CK(pwm_clk), 
            .Q(free_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i1808_1_lut (.A(n3883), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1808_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(PWMdut_m3[5]), .B(PWMdut_m3[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i17488_4_lut (.A(cnt[0]), .B(n20176), .C(cnt[2]), .D(n6), .Z(n14148)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17488_4_lut.init = 16'h0004;
    LUT4 i16778_3_lut (.A(cnt[7]), .B(n20134), .C(cnt[3]), .Z(n20176)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16778_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i16736_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n20134)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16736_4_lut.init = 16'h8000;
    LUT4 i3_4_lut (.A(n10_adj_2387), .B(PWMdut_m3[9]), .C(PWMdut_m3[8]), 
         .D(PWMdut_m3[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2316_3_lut (.A(n11440), .B(PWMdut_m3[4]), .C(PWMdut_m3[3]), 
         .Z(n10_adj_2387)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2316_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i17466_4_lut (.A(PWMdut_m3[5]), .B(n14), .C(n10_adj_2388), .D(PWMdut_m3[8]), 
         .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17466_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m3[9]), .B(PWMdut_m3[3]), .C(PWMdut_m3[4]), 
         .D(n11440), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[7]), .Z(n10_adj_2388)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_150 (.A(PWMdut_m3[2]), .B(PWMdut_m3[1]), .C(PWMdut_m3[0]), 
         .Z(n11440)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_150.init = 16'hfefe;
    CCU2D sub_1806_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m3[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18517), .S1(n3883));
    defparam sub_1806_add_2_11.INIT0 = 16'h5999;
    defparam sub_1806_add_2_11.INIT1 = 16'h0000;
    defparam sub_1806_add_2_11.INJECT1_0 = "NO";
    defparam sub_1806_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_9 (.A0(PWMdut_m3[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m3[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18516), 
          .COUT(n18517));
    defparam sub_1806_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1806_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1806_add_2_9.INJECT1_0 = "NO";
    defparam sub_1806_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_7 (.A0(PWMdut_m3[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m3[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18515), 
          .COUT(n18516));
    defparam sub_1806_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1806_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1806_add_2_7.INJECT1_0 = "NO";
    defparam sub_1806_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_5 (.A0(PWMdut_m3[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m3[4]), .C1(n9), .D1(n10), .CIN(n18514), 
          .COUT(n18515));
    defparam sub_1806_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1806_add_2_5.INIT1 = 16'h5999;
    defparam sub_1806_add_2_5.INJECT1_0 = "NO";
    defparam sub_1806_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m3[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m3[2]), .C1(n9), .D1(n10), .CIN(n18513), 
          .COUT(n18514));
    defparam sub_1806_add_2_3.INIT0 = 16'h5999;
    defparam sub_1806_add_2_3.INIT1 = 16'h5999;
    defparam sub_1806_add_2_3.INJECT1_0 = "NO";
    defparam sub_1806_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m3[0]), .C1(n9), .D1(n10), 
          .COUT(n18513));
    defparam sub_1806_add_2_1.INIT0 = 16'h0000;
    defparam sub_1806_add_2_1.INIT1 = 16'h5999;
    defparam sub_1806_add_2_1.INJECT1_0 = "NO";
    defparam sub_1806_add_2_1.INJECT1_1 = "NO";
    LUT4 i1632_3_lut_rep_390 (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .Z(n21703)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1632_3_lut_rep_390.init = 16'h1414;
    LUT4 i17524_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .D(enable_m3), .Z(n3136)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17524_2_lut_4_lut.init = 16'hebff;
    LUT4 i1602_3_lut_rep_392 (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .Z(n21705)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1602_3_lut_rep_392.init = 16'h1414;
    LUT4 i17521_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .D(enable_m3), .Z(n3100)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17521_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2105__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14148), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i0.GSR = "ENABLED";
    CCU2D cnt_2105_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18565), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2105_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2105_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2105_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2105_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18564), 
          .COUT(n18565), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2105_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2105_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2105_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2105_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18563), 
          .COUT(n18564), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2105_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2105_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2105_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2105_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18562), 
          .COUT(n18563), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2105_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2105_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2105_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2105_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18561), 
          .COUT(n18562), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2105_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2105_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2105_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2105_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18561), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2105_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2105_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2105_add_4_1.INJECT1_1 = "NO";
    FD1S3IX cnt_2105__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14148), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i1.GSR = "ENABLED";
    FD1S3IX cnt_2105__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14148), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i2.GSR = "ENABLED";
    FD1S3IX cnt_2105__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14148), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i3.GSR = "ENABLED";
    FD1S3IX cnt_2105__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14148), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i4.GSR = "ENABLED";
    FD1S3IX cnt_2105__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14148), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i5.GSR = "ENABLED";
    FD1S3IX cnt_2105__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14148), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i6.GSR = "ENABLED";
    FD1S3IX cnt_2105__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14148), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i7.GSR = "ENABLED";
    FD1S3IX cnt_2105__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14148), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i8.GSR = "ENABLED";
    FD1S3IX cnt_2105__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14148), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2105__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module HALL_U4
//

module HALL_U4 (clk_1mhz, \speed_m2[0] , hallsense_m2, rst, H_B_m2_c, 
            clkout_c_enable_272, H_A_m2_c, clkout_c_enable_341, H_C_m2_c, 
            \speed_m2[1] , \speed_m2[2] , \speed_m2[3] , \speed_m2[4] , 
            \speed_m2[5] , \speed_m2[6] , \speed_m2[7] , \speed_m2[8] , 
            \speed_m2[9] , \speed_m2[10] , \speed_m2[11] , \speed_m2[12] , 
            \speed_m2[13] , \speed_m2[14] , \speed_m2[15] , \speed_m2[16] , 
            \speed_m2[17] , \speed_m2[18] , \speed_m2[19] , GND_net, 
            n22430);
    input clk_1mhz;
    output \speed_m2[0] ;
    output [2:0]hallsense_m2;
    input rst;
    input H_B_m2_c;
    input clkout_c_enable_272;
    input H_A_m2_c;
    input clkout_c_enable_341;
    input H_C_m2_c;
    output \speed_m2[1] ;
    output \speed_m2[2] ;
    output \speed_m2[3] ;
    output \speed_m2[4] ;
    output \speed_m2[5] ;
    output \speed_m2[6] ;
    output \speed_m2[7] ;
    output \speed_m2[8] ;
    output \speed_m2[9] ;
    output \speed_m2[10] ;
    output \speed_m2[11] ;
    output \speed_m2[12] ;
    output \speed_m2[13] ;
    output \speed_m2[14] ;
    output \speed_m2[15] ;
    output \speed_m2[16] ;
    output \speed_m2[17] ;
    output \speed_m2[18] ;
    output \speed_m2[19] ;
    input GND_net;
    input n22430;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_51;
    wire [19:0]count_19__N_2067;
    
    wire stable_counting;
    wire [19:0]speedt_19__N_2047;
    
    wire hall3_lat;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4591;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21673, n21642, n4, hall2_lat, hall1_lat, hall3_old, hall1_old, 
        hall2_old, n19073, n20030, clk_1mhz_enable_186, n21, n19837, 
        n26, n22, n20164, n23, n20004, stable_counting_N_2129;
    wire [6:0]n63;
    
    wire n21691, n21647, n21650, n11466, n11464, n20180, n20178, 
        n20136, n20018, n4_adj_2386, n21675, n19928, n19803, n21638, 
        n21657, n18472, n18471, n18470, n18469, n18468, n18467, 
        n18466, n18465, n18464, n18463, n14372;
    
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2067[0]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_2047[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_19__N_2067[0]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    LUT4 i2465_2_lut_rep_329_3_lut_4_lut (.A(stable_count[3]), .B(n21673), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21642)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2465_2_lut_rep_329_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21673), .C(stable_count[0]), 
         .D(stable_count[4]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h7f8f;
    FD1P3AX hall2_lat_58 (.D(H_B_m2_c), .SP(rst), .CK(clk_1mhz), .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m2_c), .SP(clkout_c_enable_272), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m2_c), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2067[15]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2067[14]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2067[13]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2067[12]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2067[11]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2067[10]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2067[9]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2067[8]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2067[7]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2067[6]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2067[5]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2067[4]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2067[3]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2067[2]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2067[1]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2067[19]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2067[18]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2067[17]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2067[16]), .SP(clk_1mhz_enable_51), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    LUT4 i17568_4_lut (.A(n19073), .B(n20030), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_186)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17568_4_lut.init = 16'hdffd;
    FD1P3AX speed__i2 (.D(speedt_19__N_2047[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2047[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2047[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2047[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2047[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2047[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2047[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2047[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2047[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2047[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2047[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2047[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2047[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2047[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2047[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2047[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2047[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2047[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2047[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n21), .B(n19837), .C(n26), .D(n22), .Z(n19073)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i16633_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n20030)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16633_4_lut.init = 16'h7bde;
    FD1S3IX count__i1 (.D(count_19__N_2067[1]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2067[2]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2067[3]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2067[4]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2067[5]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2067[6]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2067[7]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2067[8]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2067[9]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2067[10]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2067[11]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2067[12]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2067[13]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2067[14]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2067[15]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2067[16]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2067[17]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2067[18]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2067[19]), .CK(clk_1mhz), .CD(n4591), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    LUT4 i7_2_lut (.A(count[15]), .B(n20164), .Z(n21)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i7_2_lut.init = 16'hbbbb;
    LUT4 i12_4_lut (.A(n23), .B(count[16]), .C(n20004), .D(count[1]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[17]), .B(count[4]), .C(count[18]), .D(count[6]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut (.A(count[12]), .B(count[7]), .C(count[14]), .D(count[19]), 
         .Z(n23)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2269_2_lut (.A(stable_counting), .B(stable_counting_N_2129), .Z(n4591)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2269_2_lut.init = 16'h8888;
    LUT4 i2435_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2435_1_lut.init = 16'h5555;
    LUT4 i2460_2_lut_rep_334_3_lut_4_lut (.A(stable_count[2]), .B(n21691), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21647)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2460_2_lut_rep_334_3_lut_4_lut.init = 16'h8000;
    LUT4 i2458_2_lut_rep_337_3_lut_4_lut (.A(stable_count[2]), .B(n21691), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21650)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2458_2_lut_rep_337_3_lut_4_lut.init = 16'h78f0;
    LUT4 i11517_4_lut (.A(n11466), .B(n11464), .C(stable_counting), .D(stable_counting_N_2129), 
         .Z(clk_1mhz_enable_51)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11517_4_lut.init = 16'hcaea;
    LUT4 i5_4_lut (.A(n19837), .B(n20164), .C(n20180), .D(n20178), .Z(n11466)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i5_4_lut.init = 16'h0008;
    LUT4 i16782_4_lut (.A(n20004), .B(count[15]), .C(count[14]), .D(count[18]), 
         .Z(n20180)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16782_4_lut.init = 16'hfffe;
    LUT4 i16780_4_lut (.A(count[12]), .B(n20136), .C(n20018), .D(count[19]), 
         .Z(n20178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16780_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_362 (.A(hall3_old), .B(n4_adj_2386), .C(hall3_lat), 
         .Z(n21675)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_362.init = 16'hdede;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4_adj_2386), .C(hall3_lat), 
         .D(n63[1]), .Z(n19928)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 i16738_4_lut (.A(count[17]), .B(count[7]), .C(count[6]), .D(count[1]), 
         .Z(n20136)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16738_4_lut.init = 16'hfffe;
    LUT4 i16621_2_lut (.A(count[16]), .B(count[4]), .Z(n20018)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16621_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(n21650), .B(stable_count[0]), .C(n19803), .D(n19928), 
         .Z(n11464)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2047[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2047[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2047[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2047[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2047[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2047[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2047[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2047[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2047[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_147 (.A(n21638), .B(n19928), .C(n63[2]), .D(n4), 
         .Z(stable_counting_N_2129)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_147.init = 16'h0004;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2047[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2047[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2047[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2047[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2437_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2437_2_lut.init = 16'h6666;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2047[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2047[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2047[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2047[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2047[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2047[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11466), .B(n11464), .C(count_19__N_2067[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2047[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2439_2_lut_rep_378 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21691)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2439_2_lut_rep_378.init = 16'h8888;
    LUT4 i2444_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2444_2_lut_3_lut.init = 16'h7878;
    LUT4 i2451_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2451_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2446_2_lut_rep_360_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21673)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2446_2_lut_rep_360_3_lut.init = 16'h8080;
    LUT4 i2453_2_lut_rep_344_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21657)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2453_2_lut_rep_344_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_148 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4_adj_2386)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_148.init = 16'h7bde;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18472), 
          .S0(count_19__N_2067[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18471), .COUT(n18472), .S0(count_19__N_2067[17]), .S1(count_19__N_2067[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18470), .COUT(n18471), .S0(count_19__N_2067[15]), .S1(count_19__N_2067[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18469), .COUT(n18470), .S0(count_19__N_2067[13]), .S1(count_19__N_2067[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18468), .COUT(n18469), .S0(count_19__N_2067[11]), .S1(count_19__N_2067[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    LUT4 i16607_2_lut (.A(count[11]), .B(count[5]), .Z(n20004)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16607_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(count[10]), .B(count[2]), .C(count[0]), .Z(n19837)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i16766_4_lut (.A(count[3]), .B(count[8]), .C(count[9]), .D(count[13]), 
         .Z(n20164)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16766_4_lut.init = 16'h8000;
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18467), .COUT(n18468), .S0(count_19__N_2067[9]), .S1(count_19__N_2067[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18466), 
          .COUT(n18467), .S0(count_19__N_2067[7]), .S1(count_19__N_2067[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_149 (.A(n63[3]), .B(n63[6]), .C(n21642), .D(n63[2]), 
         .Z(n19803)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_149.init = 16'hfffe;
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18465), 
          .COUT(n18466), .S0(count_19__N_2067[5]), .S1(count_19__N_2067[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_325_4_lut (.A(stable_count[5]), .B(n21647), .C(n63[6]), 
         .D(n63[3]), .Z(n21638)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_325_4_lut.init = 16'hfff6;
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18464), 
          .COUT(n18465), .S0(count_19__N_2067[3]), .S1(count_19__N_2067[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18463), 
          .COUT(n18464), .S0(count_19__N_2067[1]), .S1(count_19__N_2067[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21642), .SP(stable_counting), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21650), .SP(stable_counting), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18463), 
          .S1(count_19__N_2067[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i16752_3_lut (.A(n21675), .B(stable_counting), .C(stable_counting_N_2129), 
         .Z(n14372)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16752_3_lut.init = 16'hc8c8;
    LUT4 i2472_3_lut_4_lut (.A(stable_count[4]), .B(n21657), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2472_3_lut_4_lut.init = 16'h7f80;
    FD1P3IX stable_counting_62 (.D(n22430), .SP(clk_1mhz_enable_186), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14372), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \PID(16000000,160000000,10000000) 
//

module \PID(16000000,160000000,10000000)  (GND_net, n4466, n4465, speed_set_m3, 
            speed_set_m4, clk_N_875, n4468, n4467, n4470, n4469, 
            \subOut_24__N_1369[0] , speed_set_m2, PWMdut_m2, speed_set_m1, 
            \speed_avg_m3[12] , \speed_avg_m2[12] , \speed_avg_m3[9] , 
            \speed_avg_m2[9] , \speed_avg_m3[8] , \speed_avg_m2[8] , \speed_avg_m3[7] , 
            \speed_avg_m2[7] , \speed_avg_m3[3] , \speed_avg_m2[3] , \speed_avg_m4[19] , 
            \speed_avg_m3[19] , \speed_avg_m4[18] , \speed_avg_m3[18] , 
            \speed_avg_m4[17] , \speed_avg_m3[17] , \speed_avg_m4[16] , 
            \speed_avg_m3[16] , \speed_avg_m4[15] , \speed_avg_m3[15] , 
            \speed_avg_m4[14] , \speed_avg_m3[14] , \speed_avg_m4[13] , 
            \speed_avg_m3[13] , \speed_avg_m4[11] , \speed_avg_m3[11] , 
            \speed_avg_m4[10] , \speed_avg_m3[10] , \speed_avg_m4[6] , 
            \speed_avg_m3[6] , dir_m2, dir_m3, dir_m1, dir_m4, \speed_avg_m4[5] , 
            \speed_avg_m3[5] , \speed_avg_m4[4] , \speed_avg_m3[4] , n4472, 
            n4471, \speed_avg_m4[2] , \speed_avg_m3[2] , \speed_avg_m4[1] , 
            \speed_avg_m3[1] , \speed_avg_m4[0] , \speed_avg_m3[0] , VCC_net, 
            \speed_avg_m1[12] , \speed_avg_m1[9] , \speed_avg_m1[8] , 
            n4474, n4473, \speed_avg_m1[7] , \speed_avg_m1[3] , \speed_avg_m1[19] , 
            \speed_avg_m2[19] , \speed_avg_m1[18] , \speed_avg_m2[18] , 
            \speed_avg_m1[17] , \speed_avg_m2[17] , \speed_avg_m1[16] , 
            \speed_avg_m2[16] , \speed_avg_m1[15] , \speed_avg_m2[15] , 
            \speed_avg_m1[14] , \speed_avg_m2[14] , \speed_avg_m1[13] , 
            \speed_avg_m2[13] , \speed_avg_m1[11] , \speed_avg_m2[11] , 
            \speed_avg_m1[10] , \speed_avg_m2[10] , \speed_avg_m1[6] , 
            \speed_avg_m2[6] , \speed_avg_m1[5] , \speed_avg_m2[5] , \speed_avg_m1[4] , 
            \speed_avg_m2[4] , \speed_avg_m1[2] , \speed_avg_m2[2] , \speed_avg_m1[1] , 
            \speed_avg_m2[1] , \speed_avg_m1[0] , \speed_avg_m2[0] , n4475, 
            \subOut_24__N_1369[1] , \subOut_24__N_1369[2] , \subOut_24__N_1369[3] , 
            \subOut_24__N_1369[4] , \subOut_24__N_1369[5] , \subOut_24__N_1369[6] , 
            \subOut_24__N_1369[7] , \subOut_24__N_1369[8] , \subOut_24__N_1369[9] , 
            \subOut_24__N_1369[10] , \subOut_24__N_1369[11] , \subOut_24__N_1369[12] , 
            \subOut_24__N_1369[13] , \subOut_24__N_1369[14] , \subOut_24__N_1369[15] , 
            \subOut_24__N_1369[16] , \subOut_24__N_1369[17] , \subOut_24__N_1369[18] , 
            \subOut_24__N_1369[19] , \subOut_24__N_1369[20] , \subOut_24__N_1369[21] , 
            \subOut_24__N_1369[24] , n19942, n22435, PWMdut_m1, \speed_avg_m4[12] , 
            \speed_avg_m4[9] , \speed_avg_m4[8] , \speed_avg_m4[7] , \speed_avg_m4[3] , 
            n4479, n4481, n4480, n4483, n4482, PWMdut_m4, n4485, 
            n4484, PWMdut_m3, n4487, n4486, n4489, n4488, n4491, 
            n4490, n4493, n4492, n4495, n4494, n4497, n4496, n4499, 
            n4498, n4500, n4454, n4453, n4456, n4455, n4458, n4457, 
            n4460, n4459, n4462, n4461, n4464, n4463);
    input GND_net;
    output n4466;
    output n4465;
    input [20:0]speed_set_m3;
    input [20:0]speed_set_m4;
    input clk_N_875;
    output n4468;
    output n4467;
    output n4470;
    output n4469;
    input \subOut_24__N_1369[0] ;
    input [20:0]speed_set_m2;
    output [9:0]PWMdut_m2;
    input [20:0]speed_set_m1;
    input \speed_avg_m3[12] ;
    input \speed_avg_m2[12] ;
    input \speed_avg_m3[9] ;
    input \speed_avg_m2[9] ;
    input \speed_avg_m3[8] ;
    input \speed_avg_m2[8] ;
    input \speed_avg_m3[7] ;
    input \speed_avg_m2[7] ;
    input \speed_avg_m3[3] ;
    input \speed_avg_m2[3] ;
    input \speed_avg_m4[19] ;
    input \speed_avg_m3[19] ;
    input \speed_avg_m4[18] ;
    input \speed_avg_m3[18] ;
    input \speed_avg_m4[17] ;
    input \speed_avg_m3[17] ;
    input \speed_avg_m4[16] ;
    input \speed_avg_m3[16] ;
    input \speed_avg_m4[15] ;
    input \speed_avg_m3[15] ;
    input \speed_avg_m4[14] ;
    input \speed_avg_m3[14] ;
    input \speed_avg_m4[13] ;
    input \speed_avg_m3[13] ;
    input \speed_avg_m4[11] ;
    input \speed_avg_m3[11] ;
    input \speed_avg_m4[10] ;
    input \speed_avg_m3[10] ;
    input \speed_avg_m4[6] ;
    input \speed_avg_m3[6] ;
    output dir_m2;
    output dir_m3;
    output dir_m1;
    output dir_m4;
    input \speed_avg_m4[5] ;
    input \speed_avg_m3[5] ;
    input \speed_avg_m4[4] ;
    input \speed_avg_m3[4] ;
    output n4472;
    output n4471;
    input \speed_avg_m4[2] ;
    input \speed_avg_m3[2] ;
    input \speed_avg_m4[1] ;
    input \speed_avg_m3[1] ;
    input \speed_avg_m4[0] ;
    input \speed_avg_m3[0] ;
    input VCC_net;
    input \speed_avg_m1[12] ;
    input \speed_avg_m1[9] ;
    input \speed_avg_m1[8] ;
    output n4474;
    output n4473;
    input \speed_avg_m1[7] ;
    input \speed_avg_m1[3] ;
    input \speed_avg_m1[19] ;
    input \speed_avg_m2[19] ;
    input \speed_avg_m1[18] ;
    input \speed_avg_m2[18] ;
    input \speed_avg_m1[17] ;
    input \speed_avg_m2[17] ;
    input \speed_avg_m1[16] ;
    input \speed_avg_m2[16] ;
    input \speed_avg_m1[15] ;
    input \speed_avg_m2[15] ;
    input \speed_avg_m1[14] ;
    input \speed_avg_m2[14] ;
    input \speed_avg_m1[13] ;
    input \speed_avg_m2[13] ;
    input \speed_avg_m1[11] ;
    input \speed_avg_m2[11] ;
    input \speed_avg_m1[10] ;
    input \speed_avg_m2[10] ;
    input \speed_avg_m1[6] ;
    input \speed_avg_m2[6] ;
    input \speed_avg_m1[5] ;
    input \speed_avg_m2[5] ;
    input \speed_avg_m1[4] ;
    input \speed_avg_m2[4] ;
    input \speed_avg_m1[2] ;
    input \speed_avg_m2[2] ;
    input \speed_avg_m1[1] ;
    input \speed_avg_m2[1] ;
    input \speed_avg_m1[0] ;
    input \speed_avg_m2[0] ;
    output n4475;
    input \subOut_24__N_1369[1] ;
    input \subOut_24__N_1369[2] ;
    input \subOut_24__N_1369[3] ;
    input \subOut_24__N_1369[4] ;
    input \subOut_24__N_1369[5] ;
    input \subOut_24__N_1369[6] ;
    input \subOut_24__N_1369[7] ;
    input \subOut_24__N_1369[8] ;
    input \subOut_24__N_1369[9] ;
    input \subOut_24__N_1369[10] ;
    input \subOut_24__N_1369[11] ;
    input \subOut_24__N_1369[12] ;
    input \subOut_24__N_1369[13] ;
    input \subOut_24__N_1369[14] ;
    input \subOut_24__N_1369[15] ;
    input \subOut_24__N_1369[16] ;
    input \subOut_24__N_1369[17] ;
    input \subOut_24__N_1369[18] ;
    input \subOut_24__N_1369[19] ;
    input \subOut_24__N_1369[20] ;
    input \subOut_24__N_1369[21] ;
    input \subOut_24__N_1369[24] ;
    output n19942;
    input n22435;
    output [9:0]PWMdut_m1;
    input \speed_avg_m4[12] ;
    input \speed_avg_m4[9] ;
    input \speed_avg_m4[8] ;
    input \speed_avg_m4[7] ;
    input \speed_avg_m4[3] ;
    output n4479;
    output n4481;
    output n4480;
    output n4483;
    output n4482;
    output [9:0]PWMdut_m4;
    output n4485;
    output n4484;
    output [9:0]PWMdut_m3;
    output n4487;
    output n4486;
    output n4489;
    output n4488;
    output n4491;
    output n4490;
    output n4493;
    output n4492;
    output n4495;
    output n4494;
    output n4497;
    output n4496;
    output n4499;
    output n4498;
    output n4500;
    output n4454;
    output n4453;
    output n4456;
    output n4455;
    output n4458;
    output n4457;
    output n4460;
    output n4459;
    output n4462;
    output n4461;
    output n4464;
    output n4463;
    
    wire clk_N_875 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    wire [15:0]n1315;
    wire [9:0]n2273;
    
    wire n30;
    wire [9:0]n1451;
    
    wire n6, n22424;
    wire [28:0]intgOut1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(68[9:17])
    wire [28:0]intgOut2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(69[9:17])
    wire [28:0]n645;
    
    wire n18661;
    wire [21:0]n2353;
    
    wire n4419, n4418, n18662;
    wire [15:0]n1294;
    wire [9:0]n2261;
    
    wire n9;
    wire [9:0]n1407;
    
    wire n15564, n49;
    wire [21:0]n2593;
    
    wire n56, n22418, n21631, n18779, n18780;
    wire [28:0]backOut0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(77[9:17])
    
    wire clk_N_875_enable_72;
    wire [28:0]Out3_28__N_1174;
    wire [28:0]backOut1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(78[9:17])
    
    wire clk_N_875_enable_44, n18660, n4421, n4420;
    wire [4:0]ss;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(96[9:11])
    
    wire n21725, n21515, n18659, n4423, n4422;
    wire [28:0]multOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(88[9:16])
    wire [53:0]multOut_28__N_1411;
    
    wire n21726, n21681, n22425, n22426, n22433, n22440, n21684, 
        n21646, n21686, n21728, n21687, n19955, n21634, n16127, 
        n18417, n5440, n5442, n18418, n11474, n21635, n2545, n18416, 
        n5436, n5438, clk_N_875_enable_333;
    wire [28:0]intgOut2_28__N_1029;
    wire [28:0]intgOut3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(70[9:17])
    
    wire clk_N_875_enable_309;
    wire [28:0]intgOut3_28__N_1058;
    wire [28:0]Out0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(72[9:13])
    
    wire clk_N_875_enable_108;
    wire [28:0]Out1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(73[9:13])
    
    wire clk_N_875_enable_136;
    wire [28:0]Out2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(74[9:13])
    
    wire clk_N_875_enable_164;
    wire [28:0]Out3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(75[9:13])
    
    wire clk_N_875_enable_192;
    wire [28:0]backOut2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(79[9:17])
    
    wire clk_N_875_enable_220;
    wire [28:0]backOut3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(80[9:17])
    
    wire clk_N_875_enable_248, n19945, n16309, n42;
    wire [24:0]subOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(84[9:15])
    
    wire n21729, n21688, n5346, n3844, n1065;
    wire [28:0]addOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(92[9:15])
    wire [28:0]intgOut0_28__N_1627;
    wire [28:0]intgOut0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(67[9:17])
    
    wire clk_N_875_enable_389, n14232, n19964, n5332, n21708, n5318, 
        n5354, n22419, n14, n15, n19947, n5336, n21674, n21648;
    wire [23:0]multIn2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(87[9:16])
    
    wire n5352, n5340, n21677, n21676, n18415, n5432, n5434, clk_N_875_enable_391, 
        n18943, n30_adj_2327;
    wire [15:0]n1357;
    
    wire n14363, n22411, n5328, n5326, n5324, n14345, n5322, n5356, 
        n5350, n5348, n5342, n5358, n21731, n5344, n21721;
    wire [28:0]n585;
    
    wire n5334, n5330, n5338, n5360, subIn1_24__N_1342, n35, n21636, 
        n5392, n5400, n5368;
    wire [28:0]backOut3_28__N_1872;
    
    wire n19967, n16477, n19913, clk_N_875_enable_392, n5366, n5364, 
        n18778, n3660, n35_adj_2328, n40, n36, n4, n5320, n38, 
        n32, n34, n24, n5398, n5402, n5396, n22423;
    wire [20:0]subIn2_24__N_1534;
    
    wire n21678, n21628, n5386, n14260;
    wire [28:0]n675;
    wire [9:0]n2297;
    wire [9:0]n1539;
    
    wire n5372, n5380, n5390, n5384, n21730, n21668, n4358, n5382, 
        n5376, n34_adj_2329, n18414, n5428, n5430, n18413, n5424, 
        n5426, n18412, n5420, n5422, n18411, n5416, n5418, n18410, 
        n5412, n5414, n18406, n18407, n18408, n18409, n18405, 
        n5410, n24_adj_2330, n5374, subIn1_24__N_1533, dirout_m3_N_1947, 
        subIn1_24__N_1347, dirout_m4_N_1950;
    wire [28:0]Out0_28__N_1087;
    
    wire n18777, n18658, n4425, n4424;
    wire [28:0]Out2_28__N_1145;
    
    wire n5370, n21659, n9_adj_2331;
    wire [28:0]n555;
    
    wire n5394, n18450, n18451, n5378, n5388, n16473, n21637, 
        n4_adj_2332, n3780, n3756, n35_adj_2333, n40_adj_2334, n36_adj_2335, 
        n38_adj_2336, n32_adj_2337, n4_adj_2338, n3732, n16469, n34_adj_2339, 
        n24_adj_2340;
    wire [28:0]n121;
    
    wire n21660, mult_29s_25s_0_pp_1_2, mult_29s_25s_0_pp_2_4, mult_29s_25s_0_pp_3_6, 
        mult_29s_25s_0_pp_4_8, mult_29s_25s_0_pp_5_10, mult_29s_25s_0_pp_6_12, 
        mult_29s_25s_0_pp_7_14, mult_29s_25s_0_pp_8_16, mult_29s_25s_0_pp_9_18, 
        mult_29s_25s_0_pp_10_20, mult_29s_25s_0_pp_11_22, mult_29s_25s_0_pp_12_24, 
        mult_29s_25s_0_pp_12_25, mult_29s_25s_0_pp_12_26, mult_29s_25s_0_pp_12_27, 
        mult_29s_25s_0_pp_12_28, mult_29s_25s_0_cin_lr_2, mult_29s_25s_0_cin_lr_4, 
        mult_29s_25s_0_cin_lr_6, mult_29s_25s_0_cin_lr_8, mult_29s_25s_0_cin_lr_10, 
        mult_29s_25s_0_cin_lr_12, mult_29s_25s_0_cin_lr_14, mult_29s_25s_0_cin_lr_16, 
        mult_29s_25s_0_cin_lr_18, mult_29s_25s_0_cin_lr_20, mult_29s_25s_0_cin_lr_22, 
        co_mult_29s_25s_0_0_1, mult_29s_25s_0_pp_0_2, co_mult_29s_25s_0_0_2, 
        s_mult_29s_25s_0_0_4, mult_29s_25s_0_pp_0_4, mult_29s_25s_0_pp_0_3, 
        mult_29s_25s_0_pp_1_4, mult_29s_25s_0_pp_1_3, co_mult_29s_25s_0_0_3, 
        s_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_6, mult_29s_25s_0_pp_0_6, 
        mult_29s_25s_0_pp_0_5, mult_29s_25s_0_pp_1_6, mult_29s_25s_0_pp_1_5, 
        co_mult_29s_25s_0_0_4, s_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_8, 
        mult_29s_25s_0_pp_0_8, mult_29s_25s_0_pp_0_7, mult_29s_25s_0_pp_1_8, 
        mult_29s_25s_0_pp_1_7, co_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_10, mult_29s_25s_0_pp_0_10, mult_29s_25s_0_pp_0_9, 
        mult_29s_25s_0_pp_1_10, mult_29s_25s_0_pp_1_9, co_mult_29s_25s_0_0_6, 
        s_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_12, mult_29s_25s_0_pp_0_12, 
        mult_29s_25s_0_pp_0_11, mult_29s_25s_0_pp_1_12, mult_29s_25s_0_pp_1_11, 
        co_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_14, 
        mult_29s_25s_0_pp_0_14, mult_29s_25s_0_pp_0_13, mult_29s_25s_0_pp_1_14, 
        mult_29s_25s_0_pp_1_13, co_mult_29s_25s_0_0_8, s_mult_29s_25s_0_0_15, 
        s_mult_29s_25s_0_0_16, mult_29s_25s_0_pp_0_16, mult_29s_25s_0_pp_0_15, 
        mult_29s_25s_0_pp_1_16, mult_29s_25s_0_pp_1_15, co_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_17, s_mult_29s_25s_0_0_18, mult_29s_25s_0_pp_0_18, 
        mult_29s_25s_0_pp_0_17, mult_29s_25s_0_pp_1_18, mult_29s_25s_0_pp_1_17, 
        co_mult_29s_25s_0_0_10, s_mult_29s_25s_0_0_19, s_mult_29s_25s_0_0_20, 
        mult_29s_25s_0_pp_0_20, mult_29s_25s_0_pp_0_19, mult_29s_25s_0_pp_1_20, 
        mult_29s_25s_0_pp_1_19, co_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_21, 
        s_mult_29s_25s_0_0_22, mult_29s_25s_0_pp_0_22, mult_29s_25s_0_pp_0_21, 
        mult_29s_25s_0_pp_1_22, mult_29s_25s_0_pp_1_21, co_mult_29s_25s_0_0_12, 
        s_mult_29s_25s_0_0_23, s_mult_29s_25s_0_0_24, mult_29s_25s_0_pp_0_24, 
        mult_29s_25s_0_pp_0_23, mult_29s_25s_0_pp_1_24, mult_29s_25s_0_pp_1_23, 
        co_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_25, s_mult_29s_25s_0_0_26, 
        mult_29s_25s_0_pp_0_26, mult_29s_25s_0_pp_0_25, mult_29s_25s_0_pp_1_26, 
        mult_29s_25s_0_pp_1_25, s_mult_29s_25s_0_0_27, s_mult_29s_25s_0_0_28, 
        mult_29s_25s_0_pp_0_28, mult_29s_25s_0_pp_0_27, mult_29s_25s_0_pp_1_28, 
        mult_29s_25s_0_pp_1_27, n4_adj_2341, n3636, n16481, co_mult_29s_25s_0_1_1, 
        s_mult_29s_25s_0_1_6, mult_29s_25s_0_pp_2_6, co_mult_29s_25s_0_1_2, 
        s_mult_29s_25s_0_1_7, s_mult_29s_25s_0_1_8, mult_29s_25s_0_pp_2_8, 
        mult_29s_25s_0_pp_2_7, mult_29s_25s_0_pp_3_8, mult_29s_25s_0_pp_3_7, 
        co_mult_29s_25s_0_1_3, s_mult_29s_25s_0_1_9, s_mult_29s_25s_0_1_10, 
        mult_29s_25s_0_pp_2_10, mult_29s_25s_0_pp_2_9, mult_29s_25s_0_pp_3_10, 
        mult_29s_25s_0_pp_3_9, co_mult_29s_25s_0_1_4, s_mult_29s_25s_0_1_11, 
        s_mult_29s_25s_0_1_12, mult_29s_25s_0_pp_2_12, mult_29s_25s_0_pp_2_11, 
        mult_29s_25s_0_pp_3_12, mult_29s_25s_0_pp_3_11, co_mult_29s_25s_0_1_5, 
        s_mult_29s_25s_0_1_13, s_mult_29s_25s_0_1_14, mult_29s_25s_0_pp_2_14, 
        mult_29s_25s_0_pp_2_13, mult_29s_25s_0_pp_3_14, mult_29s_25s_0_pp_3_13, 
        co_mult_29s_25s_0_1_6, s_mult_29s_25s_0_1_15, s_mult_29s_25s_0_1_16, 
        mult_29s_25s_0_pp_2_16, mult_29s_25s_0_pp_2_15, mult_29s_25s_0_pp_3_16, 
        mult_29s_25s_0_pp_3_15, co_mult_29s_25s_0_1_7, s_mult_29s_25s_0_1_17, 
        s_mult_29s_25s_0_1_18, mult_29s_25s_0_pp_2_18, mult_29s_25s_0_pp_2_17, 
        mult_29s_25s_0_pp_3_18, mult_29s_25s_0_pp_3_17, co_mult_29s_25s_0_1_8, 
        s_mult_29s_25s_0_1_19, s_mult_29s_25s_0_1_20, mult_29s_25s_0_pp_2_20, 
        mult_29s_25s_0_pp_2_19, mult_29s_25s_0_pp_3_20, mult_29s_25s_0_pp_3_19, 
        co_mult_29s_25s_0_1_9, s_mult_29s_25s_0_1_21, s_mult_29s_25s_0_1_22, 
        mult_29s_25s_0_pp_2_22, mult_29s_25s_0_pp_2_21, mult_29s_25s_0_pp_3_22, 
        mult_29s_25s_0_pp_3_21, co_mult_29s_25s_0_1_10, s_mult_29s_25s_0_1_23, 
        s_mult_29s_25s_0_1_24, mult_29s_25s_0_pp_2_24, mult_29s_25s_0_pp_2_23, 
        mult_29s_25s_0_pp_3_24, mult_29s_25s_0_pp_3_23, co_mult_29s_25s_0_1_11, 
        s_mult_29s_25s_0_1_25, s_mult_29s_25s_0_1_26, mult_29s_25s_0_pp_2_26, 
        mult_29s_25s_0_pp_2_25, mult_29s_25s_0_pp_3_26, mult_29s_25s_0_pp_3_25, 
        s_mult_29s_25s_0_1_27, s_mult_29s_25s_0_1_28, mult_29s_25s_0_pp_2_28, 
        mult_29s_25s_0_pp_2_27, mult_29s_25s_0_pp_3_28, mult_29s_25s_0_pp_3_27, 
        co_mult_29s_25s_0_2_1, s_mult_29s_25s_0_2_10, mult_29s_25s_0_pp_4_10, 
        co_mult_29s_25s_0_2_2, s_mult_29s_25s_0_2_12, s_mult_29s_25s_0_2_11, 
        mult_29s_25s_0_pp_4_12, mult_29s_25s_0_pp_4_11, mult_29s_25s_0_pp_5_12, 
        mult_29s_25s_0_pp_5_11, co_mult_29s_25s_0_2_3, s_mult_29s_25s_0_2_13, 
        s_mult_29s_25s_0_2_14, mult_29s_25s_0_pp_4_14, mult_29s_25s_0_pp_4_13, 
        mult_29s_25s_0_pp_5_14, mult_29s_25s_0_pp_5_13, co_mult_29s_25s_0_2_4, 
        s_mult_29s_25s_0_2_15, s_mult_29s_25s_0_2_16, mult_29s_25s_0_pp_4_16, 
        mult_29s_25s_0_pp_4_15, mult_29s_25s_0_pp_5_16, mult_29s_25s_0_pp_5_15, 
        co_mult_29s_25s_0_2_5, s_mult_29s_25s_0_2_17, s_mult_29s_25s_0_2_18, 
        mult_29s_25s_0_pp_4_18, mult_29s_25s_0_pp_4_17, mult_29s_25s_0_pp_5_18, 
        mult_29s_25s_0_pp_5_17, co_mult_29s_25s_0_2_6, s_mult_29s_25s_0_2_19, 
        s_mult_29s_25s_0_2_20, mult_29s_25s_0_pp_4_20, mult_29s_25s_0_pp_4_19, 
        mult_29s_25s_0_pp_5_20, mult_29s_25s_0_pp_5_19, co_mult_29s_25s_0_2_7, 
        s_mult_29s_25s_0_2_21, s_mult_29s_25s_0_2_22, mult_29s_25s_0_pp_4_22, 
        mult_29s_25s_0_pp_4_21, mult_29s_25s_0_pp_5_22, mult_29s_25s_0_pp_5_21, 
        co_mult_29s_25s_0_2_8, s_mult_29s_25s_0_2_23, s_mult_29s_25s_0_2_24, 
        mult_29s_25s_0_pp_4_24, mult_29s_25s_0_pp_4_23, mult_29s_25s_0_pp_5_24, 
        mult_29s_25s_0_pp_5_23, co_mult_29s_25s_0_2_9, s_mult_29s_25s_0_2_25, 
        s_mult_29s_25s_0_2_26, mult_29s_25s_0_pp_4_26, mult_29s_25s_0_pp_4_25, 
        mult_29s_25s_0_pp_5_26, mult_29s_25s_0_pp_5_25, s_mult_29s_25s_0_2_27, 
        s_mult_29s_25s_0_2_28, mult_29s_25s_0_pp_4_28, mult_29s_25s_0_pp_4_27, 
        mult_29s_25s_0_pp_5_28, mult_29s_25s_0_pp_5_27, n3684, co_mult_29s_25s_0_3_1, 
        s_mult_29s_25s_0_3_14, mult_29s_25s_0_pp_6_14, co_mult_29s_25s_0_3_2, 
        s_mult_29s_25s_0_3_15, s_mult_29s_25s_0_3_16, mult_29s_25s_0_pp_6_16, 
        mult_29s_25s_0_pp_6_15, mult_29s_25s_0_pp_7_16, mult_29s_25s_0_pp_7_15, 
        co_mult_29s_25s_0_3_3, s_mult_29s_25s_0_3_17, s_mult_29s_25s_0_3_18, 
        mult_29s_25s_0_pp_6_18, mult_29s_25s_0_pp_6_17, mult_29s_25s_0_pp_7_18, 
        mult_29s_25s_0_pp_7_17, co_mult_29s_25s_0_3_4, s_mult_29s_25s_0_3_19, 
        s_mult_29s_25s_0_3_20, mult_29s_25s_0_pp_6_20, mult_29s_25s_0_pp_6_19, 
        mult_29s_25s_0_pp_7_20, mult_29s_25s_0_pp_7_19, co_mult_29s_25s_0_3_5, 
        s_mult_29s_25s_0_3_21, s_mult_29s_25s_0_3_22, mult_29s_25s_0_pp_6_22, 
        mult_29s_25s_0_pp_6_21, mult_29s_25s_0_pp_7_22, mult_29s_25s_0_pp_7_21, 
        co_mult_29s_25s_0_3_6, s_mult_29s_25s_0_3_23, s_mult_29s_25s_0_3_24, 
        mult_29s_25s_0_pp_6_24, mult_29s_25s_0_pp_6_23, mult_29s_25s_0_pp_7_24, 
        mult_29s_25s_0_pp_7_23, co_mult_29s_25s_0_3_7, s_mult_29s_25s_0_3_25, 
        s_mult_29s_25s_0_3_26, mult_29s_25s_0_pp_6_26, mult_29s_25s_0_pp_6_25, 
        mult_29s_25s_0_pp_7_26, mult_29s_25s_0_pp_7_25, s_mult_29s_25s_0_3_27, 
        s_mult_29s_25s_0_3_28, mult_29s_25s_0_pp_6_28, mult_29s_25s_0_pp_6_27, 
        mult_29s_25s_0_pp_7_28, mult_29s_25s_0_pp_7_27, co_mult_29s_25s_0_4_1, 
        s_mult_29s_25s_0_4_18, mult_29s_25s_0_pp_8_18, co_mult_29s_25s_0_4_2, 
        s_mult_29s_25s_0_4_20, s_mult_29s_25s_0_4_19, mult_29s_25s_0_pp_8_20, 
        mult_29s_25s_0_pp_8_19, mult_29s_25s_0_pp_9_20, mult_29s_25s_0_pp_9_19, 
        co_mult_29s_25s_0_4_3, s_mult_29s_25s_0_4_21, s_mult_29s_25s_0_4_22, 
        mult_29s_25s_0_pp_8_22, mult_29s_25s_0_pp_8_21, mult_29s_25s_0_pp_9_22, 
        mult_29s_25s_0_pp_9_21, co_mult_29s_25s_0_4_4, s_mult_29s_25s_0_4_23, 
        s_mult_29s_25s_0_4_24, mult_29s_25s_0_pp_8_24, mult_29s_25s_0_pp_8_23, 
        mult_29s_25s_0_pp_9_24, mult_29s_25s_0_pp_9_23, co_mult_29s_25s_0_4_5, 
        s_mult_29s_25s_0_4_25, s_mult_29s_25s_0_4_26, mult_29s_25s_0_pp_8_26, 
        mult_29s_25s_0_pp_8_25, mult_29s_25s_0_pp_9_26, mult_29s_25s_0_pp_9_25, 
        s_mult_29s_25s_0_4_27, s_mult_29s_25s_0_4_28, mult_29s_25s_0_pp_8_28, 
        mult_29s_25s_0_pp_8_27, mult_29s_25s_0_pp_9_28, mult_29s_25s_0_pp_9_27, 
        co_mult_29s_25s_0_5_1, s_mult_29s_25s_0_5_22, mult_29s_25s_0_pp_10_22, 
        co_mult_29s_25s_0_5_2, s_mult_29s_25s_0_5_23, s_mult_29s_25s_0_5_24, 
        mult_29s_25s_0_pp_10_24, mult_29s_25s_0_pp_10_23, mult_29s_25s_0_pp_11_24, 
        mult_29s_25s_0_pp_11_23, co_mult_29s_25s_0_5_3, s_mult_29s_25s_0_5_25, 
        s_mult_29s_25s_0_5_26, mult_29s_25s_0_pp_10_26, mult_29s_25s_0_pp_10_25, 
        mult_29s_25s_0_pp_11_26, mult_29s_25s_0_pp_11_25, s_mult_29s_25s_0_5_27, 
        s_mult_29s_25s_0_5_28, mult_29s_25s_0_pp_10_28, mult_29s_25s_0_pp_10_27, 
        mult_29s_25s_0_pp_11_28, mult_29s_25s_0_pp_11_27, co_mult_29s_25s_0_6_1, 
        s_mult_29s_25s_0_6_24, co_mult_29s_25s_0_6_2, s_mult_29s_25s_0_6_25, 
        s_mult_29s_25s_0_6_26, s_mult_29s_25s_0_6_27, s_mult_29s_25s_0_6_28, 
        co_mult_29s_25s_0_7_1, co_mult_29s_25s_0_7_2, mult_29s_25s_0_pp_2_5, 
        co_mult_29s_25s_0_7_3, s_mult_29s_25s_0_7_8, co_mult_29s_25s_0_7_4, 
        s_mult_29s_25s_0_7_9, s_mult_29s_25s_0_7_10, co_mult_29s_25s_0_7_5, 
        s_mult_29s_25s_0_7_11, s_mult_29s_25s_0_7_12, co_mult_29s_25s_0_7_6, 
        s_mult_29s_25s_0_7_13, s_mult_29s_25s_0_7_14, co_mult_29s_25s_0_7_7, 
        s_mult_29s_25s_0_7_15, s_mult_29s_25s_0_7_16, co_mult_29s_25s_0_7_8, 
        s_mult_29s_25s_0_7_17, s_mult_29s_25s_0_7_18, co_mult_29s_25s_0_7_9, 
        s_mult_29s_25s_0_7_19, s_mult_29s_25s_0_7_20, co_mult_29s_25s_0_7_10, 
        s_mult_29s_25s_0_7_21, s_mult_29s_25s_0_7_22, co_mult_29s_25s_0_7_11, 
        s_mult_29s_25s_0_7_23, s_mult_29s_25s_0_7_24, co_mult_29s_25s_0_7_12, 
        s_mult_29s_25s_0_7_25, s_mult_29s_25s_0_7_26, s_mult_29s_25s_0_7_27, 
        s_mult_29s_25s_0_7_28, co_mult_29s_25s_0_8_1, s_mult_29s_25s_0_8_12, 
        co_mult_29s_25s_0_8_2, s_mult_29s_25s_0_8_13, s_mult_29s_25s_0_8_14, 
        mult_29s_25s_0_pp_6_13, co_mult_29s_25s_0_8_3, s_mult_29s_25s_0_8_15, 
        s_mult_29s_25s_0_8_16, co_mult_29s_25s_0_8_4, s_mult_29s_25s_0_8_17, 
        s_mult_29s_25s_0_8_18, co_mult_29s_25s_0_8_5, s_mult_29s_25s_0_8_19, 
        s_mult_29s_25s_0_8_20, co_mult_29s_25s_0_8_6, s_mult_29s_25s_0_8_21, 
        s_mult_29s_25s_0_8_22, co_mult_29s_25s_0_8_7, s_mult_29s_25s_0_8_23, 
        s_mult_29s_25s_0_8_24, co_mult_29s_25s_0_8_8, s_mult_29s_25s_0_8_25, 
        s_mult_29s_25s_0_8_26, s_mult_29s_25s_0_8_27, s_mult_29s_25s_0_8_28, 
        n16337, co_mult_29s_25s_0_9_1, s_mult_29s_25s_0_9_20, co_mult_29s_25s_0_9_2, 
        s_mult_29s_25s_0_9_21, s_mult_29s_25s_0_9_22, mult_29s_25s_0_pp_10_21, 
        co_mult_29s_25s_0_9_3, s_mult_29s_25s_0_9_24, s_mult_29s_25s_0_9_23, 
        co_mult_29s_25s_0_9_4, s_mult_29s_25s_0_9_25, s_mult_29s_25s_0_9_26, 
        s_mult_29s_25s_0_9_27, s_mult_29s_25s_0_9_28;
    wire [20:0]subIn2_24__N_1348;
    
    wire co_mult_29s_25s_0_10_1, co_mult_29s_25s_0_10_2, mult_29s_25s_0_pp_4_9, 
        co_mult_29s_25s_0_10_3, co_mult_29s_25s_0_10_4, co_mult_29s_25s_0_10_5, 
        s_mult_29s_25s_0_10_16, co_mult_29s_25s_0_10_6, s_mult_29s_25s_0_10_17, 
        s_mult_29s_25s_0_10_18, co_mult_29s_25s_0_10_7, s_mult_29s_25s_0_10_19, 
        s_mult_29s_25s_0_10_20, co_mult_29s_25s_0_10_8, s_mult_29s_25s_0_10_21, 
        s_mult_29s_25s_0_10_22, co_mult_29s_25s_0_10_9, s_mult_29s_25s_0_10_23, 
        s_mult_29s_25s_0_10_24, co_mult_29s_25s_0_10_10, s_mult_29s_25s_0_10_25, 
        s_mult_29s_25s_0_10_26, s_mult_29s_25s_0_10_27, s_mult_29s_25s_0_10_28, 
        n18657, n4427, n4426, co_mult_29s_25s_0_11_1, s_mult_29s_25s_0_11_24, 
        co_mult_29s_25s_0_11_2, s_mult_29s_25s_0_11_25, s_mult_29s_25s_0_11_26, 
        s_mult_29s_25s_0_11_27, s_mult_29s_25s_0_11_28, co_t_mult_29s_25s_0_12_1, 
        co_t_mult_29s_25s_0_12_2, mult_29s_25s_0_pp_8_17, co_t_mult_29s_25s_0_12_3, 
        co_t_mult_29s_25s_0_12_4, co_t_mult_29s_25s_0_12_5, co_t_mult_29s_25s_0_12_6, 
        mult_29s_25s_0_cin_lr_0, mco, mco_1, mco_2, mco_3, mco_4, 
        mco_5, mco_6, mco_7, mco_8, mco_9, mco_10, mco_11, mco_12, 
        mco_14, mco_15, mco_16, mco_17, mco_18, mco_19, mco_20, 
        mco_21, mco_22, mco_23, mco_24, mco_25, mco_28, mco_29, 
        mco_30, mco_31, mco_32, mco_33, mco_34, mco_35, mco_36, 
        mco_37, mco_38, mco_42, mco_43, mco_44, mco_45, mco_46, 
        mco_47, mco_48, mco_49, mco_50, mco_51, mco_56, mco_57, 
        mco_58, mco_59, mco_60, mco_61, mco_62, mco_63, mco_64, 
        mco_70, mco_71, mco_72, mco_73, mco_74, mco_75, mco_76, 
        mco_77, n5821, mco_84, mco_85, mco_86, mco_87, mco_88, 
        mco_89, mco_90, mco_98, mco_99, mco_100, mco_101, mco_102, 
        mco_103, mco_112, mco_113, mco_114, mco_115, mco_116, mco_126, 
        mco_127, mco_128, mco_129, mco_140, mco_141, mco_142, n22420, 
        n22421, mco_154, mco_155, n21630, n5518, n19907, n21697, 
        n20645, n20372, n5805, n5807, n5809, n5811, n5813, n5815, 
        n5817, n5819, n4428, n18656, n5823, n18655, n18654, n18653, 
        n16073, n18652, n18651, n5825, n18768, n18767, n18766, 
        n18650, n18765, n5827, n21666, n21723, n5829, n18649, 
        n5831, n18764, n5833, n18763, n18762, n18648, n18647, 
        n18761, n18760, n18759, n18646, n3612, n18645, n18644, 
        n18758, n5835, n5837, n5839, n5841, n5845, n18643, n18757, 
        n16131, n35_adj_2342, n40_adj_2343, n36_adj_2344, n38_adj_2345, 
        n32_adj_2346, n34_adj_2347, n24_adj_2348, n18756, n18755, 
        n18642, n4_adj_2349, n21633, n21632, n14_adj_2350, n10, 
        n18960, n6_adj_2351, n18961, n14_adj_2352, n10_adj_2353, n18945, 
        n6_adj_2354, n18946, n14_adj_2355, n10_adj_2356, n18920, n6_adj_2357, 
        n18921, n16283, n14336, n21658, n9_adj_2358, n8, n10_adj_2359, 
        n8_adj_2360, n4_adj_2361, n18641, n18640, n18639, n18638, 
        n18637, n18636, n18635, n21694, n18449, n18634, n18633, 
        n18427, n18428, n21698, n18426, n14237, n18632, n14265, 
        n18631, n18630, n18629, n18736, n18735, n9_adj_2362, n7, 
        n10_adj_2363, n18734, n8_adj_2364, n4_adj_2365, n18628, n18627, 
        n18626, n14313, n14289, n20659, n18625, n18624, n18733, 
        n18732, n18623, n18448, n18622, n18731, n18730, n18729, 
        n18728, n18727, n18621, n18447, n22427, n18726, n18446, 
        n18445, n18425, n18620, n18619, n18725, n18618, n18617, 
        n18724, n18723, n18722, n18616, n18615, n18614, n18613, 
        n18721, n18720, n18612, n18611, n18610, n18609, n18719, 
        n18718, n18717, n18716, n18715, n18714, n18713, n18712, 
        n18711, n18710, n18444;
    wire [15:0]n1336;
    
    wire n18443, n18442, n18424, n18423, n18441, n18812, n3708, 
        n18709, n18708, n18507, n18707, n18706, n18811, n18810, 
        n18506, n18705, n18704, n18703, n18809, n18808, n18702, 
        n18701, n18700, n18807, n18806, n18589;
    wire [28:0]addIn2_28__N_1440;
    
    wire n18505, n18588, n18587, n18699, n18504, n18805, n18698, 
        n18586, n18585, n18697, n18804, n18440, n18503, n18584, 
        n18439, n18583, n18696, n18438, n18803, n18802, n18582, 
        n18422, n18581, n18801, n18580, n18800, n18799, n18502;
    wire [9:0]n2285;
    
    wire n18501, n18579, n18578, n18577, n18798, n18797, n18500, 
        n14_adj_2366, n10_adj_2367, n18892, n18499, n18576, n18687, 
        n5450, n18686, n5448, n5446, n5444, n6_adj_2368, n18893, 
        n18685, n18684, n18796, n18795, n14340, n5519, n5806, 
        n5808, n5810, n5812, n5814, n5816;
    wire [20:0]n367;
    
    wire n5818, n18683, n18682, n5820, n18498, n18681, n5822, 
        n18680, n5824, n18421, n5826, n5828, n5830, n5832, n5834, 
        n18497, n18496, n18495, n18494, n18437, n18679, n8_adj_2369, 
        n5846, n5836, n5838, n5840, n5842;
    wire [28:0]n615;
    wire [28:0]addIn2_28__N_1569;
    
    wire n20384, n18493, n18678, n4409, n18677, n4411, n4410, 
        n19337, n19331, n19325, n18676, n4413, n4412;
    wire [9:0]n1495;
    
    wire n18675, n4415, n4414, n14354, n19319, n19313, n19307, 
        n18674, n4417, n4416, n18673, n18672, n9_adj_2370, n7_adj_2371, 
        n10_adj_2372, n8_adj_2373, n4_adj_2374, n18671, n9_adj_2375, 
        n18436, n9_adj_2376, n8_adj_2377, n10_adj_2378, n8_adj_2379, 
        n4_adj_2380, n35_adj_2381, n40_adj_2382, n36_adj_2383, n21737, 
        n21736, n38_adj_2384, n32_adj_2385, n18435, n18670, n18669, 
        n18667, n18434, n18420, n18419, n18433, n18432, n18431, 
        n18430, n18666, n18665, n18429, n18664, n18784, n18663, 
        n18783, n18782, n18452, n18781;
    
    LUT4 i1_3_lut (.A(n1315[15]), .B(n2273[6]), .C(n30), .Z(n1451[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut.init = 16'h8a8a;
    LUT4 mux_138_i29_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[28]), 
         .D(intgOut2[28]), .Z(n645[28])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i29_3_lut_4_lut.init = 16'hfe10;
    CCU2D sub_16_rep_3_add_2_11 (.A0(n2353[9]), .B0(n4419), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[10]), .B1(n4418), .C1(GND_net), .D1(GND_net), 
          .CIN(n18661), .COUT(n18662), .S0(n4466), .S1(n4465));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_11.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_11.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_11.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_42 (.A(n1294[15]), .B(n2261[9]), .C(n9), .Z(n1407[9])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_42.init = 16'h8a8a;
    LUT4 mux_1253_i4_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[3]), 
         .D(speed_set_m4[3]), .Z(n2593[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1253_i11_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[10]), 
         .D(speed_set_m4[10]), .Z(n2593[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_adj_43 (.A(n1294[15]), .B(n2261[8]), .C(n9), .Z(n1407[8])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_43.init = 16'h8a8a;
    LUT4 i1_2_lut_rep_318_3_lut_4_lut (.A(n15564), .B(n49), .C(n56), .D(n22418), 
         .Z(n21631)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i1_2_lut_rep_318_3_lut_4_lut.init = 16'heee0;
    LUT4 i1_3_lut_adj_44 (.A(n1294[15]), .B(n2261[7]), .C(n9), .Z(n1407[7])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_44.init = 16'h8a8a;
    LUT4 mux_1253_i5_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[4]), 
         .D(speed_set_m4[4]), .Z(n2593[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i5_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15369_7 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18779), .COUT(n18780));
    defparam add_15369_7.INIT0 = 16'h0aaa;
    defparam add_15369_7.INIT1 = 16'hf555;
    defparam add_15369_7.INJECT1_0 = "NO";
    defparam add_15369_7.INJECT1_1 = "NO";
    FD1P3AX backOut0_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_adj_45 (.A(n1294[15]), .B(n2261[6]), .C(n9), .Z(n1407[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_45.init = 16'h8a8a;
    LUT4 mux_1253_i6_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[5]), 
         .D(speed_set_m4[5]), .Z(n2593[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i5_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[4]), 
         .D(intgOut2[4]), .Z(n645[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i5_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_adj_46 (.A(n1294[15]), .B(n2261[5]), .C(n9), .Z(n1407[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_46.init = 16'h8a8a;
    FD1P3AX backOut1_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_adj_47 (.A(n1294[15]), .B(n2261[3]), .C(n9), .Z(n1407[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_47.init = 16'h8a8a;
    LUT4 mux_138_i22_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[21]), 
         .D(intgOut2[21]), .Z(n645[21])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i22_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i17_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[16]), 
         .D(intgOut2[16]), .Z(n645[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i17_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i14_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[13]), 
         .D(intgOut2[13]), .Z(n645[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i14_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1253_i15_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[14]), 
         .D(speed_set_m4[14]), .Z(n2593[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i20_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[19]), 
         .D(intgOut2[19]), .Z(n645[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i20_3_lut_4_lut.init = 16'hfe10;
    CCU2D sub_16_rep_3_add_2_9 (.A0(n2353[7]), .B0(n4421), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[8]), .B1(n4420), .C1(GND_net), .D1(GND_net), 
          .CIN(n18660), .COUT(n18661), .S0(n4468), .S1(n4467));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_9.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_9.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_412 (.A(ss[0]), .B(ss[3]), .Z(n21725)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_412.init = 16'h8888;
    LUT4 ss_2__bdd_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), .D(ss[2]), 
         .Z(n21515)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam ss_2__bdd_3_lut_4_lut.init = 16'h0800;
    CCU2D sub_16_rep_3_add_2_7 (.A0(n2353[5]), .B0(n4423), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[6]), .B1(n4422), .C1(GND_net), .D1(GND_net), 
          .CIN(n18659), .COUT(n18660), .S0(n4470), .S1(n4469));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_7.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_7.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_7.INJECT1_1 = "NO";
    LUT4 mux_138_i23_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[22]), 
         .D(intgOut2[22]), .Z(n645[22])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i23_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i26_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[25]), 
         .D(intgOut2[25]), .Z(n645[25])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i26_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i4_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[3]), 
         .D(intgOut2[3]), .Z(n645[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i28_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[27]), 
         .D(intgOut2[27]), .Z(n645[27])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i28_3_lut_4_lut.init = 16'hfe10;
    FD1S3AX multOut_i0 (.D(multOut_28__N_1411[0]), .CK(clk_N_875), .Q(multOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_413 (.A(ss[1]), .B(ss[2]), .Z(n21726)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_413.init = 16'h2222;
    LUT4 mux_138_i6_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[5]), 
         .D(intgOut2[5]), .Z(n645[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1253_i1_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[0]), 
         .D(speed_set_m4[0]), .Z(n2593[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i7_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[6]), 
         .D(intgOut2[6]), .Z(n645[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 i2_3_lut_rep_335_4_lut_else_3_lut (.A(n21681), .B(ss[3]), .C(n22425), 
         .D(ss[1]), .Z(n22426)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C (D))+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(174[9:17])
    defparam i2_3_lut_rep_335_4_lut_else_3_lut.init = 16'hf3aa;
    LUT4 i1_2_lut_rep_371_3_lut (.A(n22433), .B(n22440), .C(ss[3]), .Z(n21684)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_371_3_lut.init = 16'hefef;
    LUT4 i17583_2_lut_rep_333_2_lut_3_lut_4_lut (.A(n22433), .B(n22440), 
         .C(n6), .D(ss[3]), .Z(n21646)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i17583_2_lut_rep_333_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_373_3_lut (.A(n22433), .B(n22440), .C(ss[3]), .Z(n21686)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_373_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_415 (.A(ss[0]), .B(ss[3]), .Z(n21728)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_415.init = 16'hbbbb;
    LUT4 i2_2_lut_rep_374_3_lut (.A(ss[0]), .B(ss[3]), .C(n22433), .Z(n21687)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_2_lut_rep_374_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n19955)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i52_2_lut_rep_321 (.A(n15564), .B(n49), .Z(n21634)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(138[23] 139[51])
    defparam i52_2_lut_rep_321.init = 16'h4444;
    LUT4 mux_138_i11_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[10]), 
         .D(intgOut2[10]), .Z(n645[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13562_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), .D(ss[2]), 
         .Z(n16127)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13562_2_lut_3_lut_4_lut.init = 16'hfffb;
    CCU2D add_1188_17 (.A0(n5440), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5442), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18417), 
          .COUT(n18418), .S0(n2353[15]), .S1(n2353[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_17.INIT0 = 16'hf555;
    defparam add_1188_17.INIT1 = 16'hf555;
    defparam add_1188_17.INJECT1_0 = "NO";
    defparam add_1188_17.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(n15564), .B(n49), .C(n11474), .D(n21635), 
         .Z(n2545)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(138[23] 139[51])
    defparam i1_3_lut_4_lut.init = 16'hf040;
    LUT4 mux_138_i12_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[11]), 
         .D(intgOut2[11]), .Z(n645[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i12_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1188_15 (.A0(n5436), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5438), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18416), 
          .COUT(n18417), .S0(n2353[13]), .S1(n2353[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_15.INIT0 = 16'hf555;
    defparam add_1188_15.INIT1 = 16'hf555;
    defparam add_1188_15.INJECT1_0 = "NO";
    defparam add_1188_15.INJECT1_1 = "NO";
    LUT4 mux_138_i13_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[12]), 
         .D(intgOut2[12]), .Z(n645[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i13_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX intgOut2_i0 (.D(intgOut2_28__N_1029[0]), .SP(clk_N_875_enable_333), 
            .CK(clk_N_875), .Q(intgOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i0.GSR = "ENABLED";
    FD1P3AX intgOut3_i0 (.D(intgOut3_28__N_1058[0]), .SP(clk_N_875_enable_309), 
            .CK(clk_N_875), .Q(intgOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i0.GSR = "ENABLED";
    FD1P3AX Out0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i0.GSR = "ENABLED";
    FD1P3AX Out1_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i0.GSR = "ENABLED";
    FD1P3AX Out2_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i0.GSR = "ENABLED";
    FD1P3AX Out3_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i0.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i0.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .D(ss[1]), 
         .Z(n19945)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_322 (.A(n16309), .B(n42), .Z(n21635)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam i1_2_lut_rep_322.init = 16'h4444;
    FD1S3AX subOut_i0 (.D(\subOut_24__N_1369[0] ), .CK(clk_N_875), .Q(subOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i0.GSR = "ENABLED";
    LUT4 i13026_2_lut_rep_416 (.A(n22440), .B(ss[3]), .Z(n21729)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13026_2_lut_rep_416.init = 16'heeee;
    LUT4 mux_138_i16_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[15]), 
         .D(intgOut2[15]), .Z(n645[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i19_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[18]), 
         .D(intgOut2[18]), .Z(n645[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i19_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i21_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[20]), 
         .D(intgOut2[20]), .Z(n645[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i24_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[23]), 
         .D(intgOut2[23]), .Z(n645[23])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i24_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i25_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[24]), 
         .D(intgOut2[24]), .Z(n645[24])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_rep_375_3_lut_4_lut (.A(n22440), .B(ss[3]), .C(ss[1]), 
         .D(ss[0]), .Z(n21688)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_rep_375_3_lut_4_lut.init = 16'h0110;
    LUT4 mux_1198_i14_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[13]), 
         .D(speed_set_m3[13]), .Z(n5346)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i2_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[1]), 
         .D(intgOut2[1]), .Z(n645[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i2_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i3_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[2]), 
         .D(intgOut2[2]), .Z(n645[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i27_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[26]), 
         .D(intgOut2[26]), .Z(n645[26])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i27_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i8_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[7]), 
         .D(intgOut2[7]), .Z(n645[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3111_3_lut (.A(n3844), .B(n1065), .C(addOut[28]), .Z(intgOut0_28__N_1627[28])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3111_3_lut.init = 16'h3232;
    FD1P3IX intgOut0_i0 (.D(addOut[0]), .SP(clk_N_875_enable_389), .CD(n14232), 
            .CK(clk_N_875), .Q(intgOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i0.GSR = "ENABLED";
    LUT4 mux_138_i1_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[0]), 
         .D(intgOut2[0]), .Z(n645[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut (.A(n22440), .B(ss[1]), .Z(n19964)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 mux_1198_i7_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[6]), 
         .D(speed_set_m3[6]), .Z(n5332)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i7_3_lut_4_lut.init = 16'hfb40;
    FD1S3IX ss_i0 (.D(n21708), .CK(clk_N_875), .CD(ss[4]), .Q(ss[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i0.GSR = "ENABLED";
    LUT4 mux_1198_i1_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[0]), 
         .D(speed_set_m3[0]), .Z(n5318)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i18_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[17]), 
         .D(speed_set_m3[17]), .Z(n5354)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i18_3_lut_4_lut.init = 16'hfb40;
    FD1S3IX ss_i1 (.D(n22419), .CK(clk_N_875), .CD(ss[4]), .Q(ss[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i1.GSR = "ENABLED";
    FD1S3IX ss_i2 (.D(n14), .CK(clk_N_875), .CD(ss[4]), .Q(ss[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i2.GSR = "ENABLED";
    FD1S3IX ss_i3 (.D(n15), .CK(clk_N_875), .CD(ss[4]), .Q(ss[3]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i3.GSR = "ENABLED";
    FD1S3AY ss_i4 (.D(n19947), .CK(clk_N_875), .Q(ss[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i4.GSR = "ENABLED";
    LUT4 mux_1198_i9_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[8]), 
         .D(speed_set_m3[8]), .Z(n5336)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3109_3_lut (.A(n3844), .B(n1065), .C(addOut[27]), .Z(intgOut0_28__N_1627[27])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3109_3_lut.init = 16'h3232;
    LUT4 i3107_3_lut (.A(n3844), .B(n1065), .C(addOut[26]), .Z(intgOut0_28__N_1627[26])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3107_3_lut.init = 16'h3232;
    LUT4 i3105_3_lut (.A(n3844), .B(n1065), .C(addOut[25]), .Z(intgOut0_28__N_1627[25])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3105_3_lut.init = 16'h3232;
    LUT4 i17544_2_lut_3_lut_4_lut_4_lut (.A(n21674), .B(n21648), .C(n21681), 
         .D(n6), .Z(multIn2[2])) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i17544_2_lut_3_lut_4_lut_4_lut.init = 16'h1115;
    LUT4 mux_1198_i17_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[16]), 
         .D(speed_set_m3[16]), .Z(n5352)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i11_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[10]), 
         .D(speed_set_m3[10]), .Z(n5340)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_4_lut (.A(n21677), .B(n22440), .C(n21676), .D(ss[3]), 
         .Z(clk_N_875_enable_192)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam i1_4_lut_4_lut.init = 16'hb888;
    LUT4 i1_4_lut_4_lut_adj_48 (.A(n21677), .B(n22440), .C(n19955), .D(ss[1]), 
         .Z(clk_N_875_enable_164)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(B+(C+!(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_48.init = 16'h8b88;
    LUT4 i1_4_lut_4_lut_adj_49 (.A(n21677), .B(n22440), .C(n19955), .D(ss[1]), 
         .Z(clk_N_875_enable_108)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+(C+(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_49.init = 16'h888b;
    CCU2D add_1188_13 (.A0(n5432), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5434), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18415), 
          .COUT(n18416), .S0(n2353[11]), .S1(n2353[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_13.INIT0 = 16'hf555;
    defparam add_1188_13.INIT1 = 16'hf555;
    defparam add_1188_13.INJECT1_0 = "NO";
    defparam add_1188_13.INJECT1_1 = "NO";
    LUT4 i3103_3_lut (.A(n3844), .B(n1065), .C(addOut[24]), .Z(intgOut0_28__N_1627[24])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3103_3_lut.init = 16'h3232;
    LUT4 i3101_3_lut (.A(n3844), .B(n1065), .C(addOut[23]), .Z(intgOut0_28__N_1627[23])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3101_3_lut.init = 16'h3232;
    LUT4 i3099_3_lut (.A(n3844), .B(n1065), .C(addOut[22]), .Z(intgOut0_28__N_1627[22])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3099_3_lut.init = 16'h3232;
    LUT4 i11778_4_lut (.A(clk_N_875_enable_391), .B(n18943), .C(n30_adj_2327), 
         .D(n1357[15]), .Z(n14363)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11778_4_lut.init = 16'h8aaa;
    LUT4 ss_3__bdd_4_lut (.A(ss[3]), .B(n22433), .C(ss[0]), .D(ss[1]), 
         .Z(n22411)) /* synthesis lut_function=(A (C+(D))+!A !(B (C (D)))) */ ;
    defparam ss_3__bdd_4_lut.init = 16'hbff5;
    LUT4 mux_1198_i5_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[4]), 
         .D(speed_set_m3[4]), .Z(n5328)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3097_3_lut (.A(n3844), .B(n1065), .C(addOut[21]), .Z(intgOut0_28__N_1627[21])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3097_3_lut.init = 16'h3232;
    LUT4 mux_1198_i4_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[3]), 
         .D(speed_set_m3[3]), .Z(n5326)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i3_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[2]), 
         .D(speed_set_m3[2]), .Z(n5324)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i3_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX dutyout_m2_i0_i0 (.D(n2273[0]), .SP(clk_N_875_enable_391), .CD(n14345), 
            .CK(clk_N_875), .Q(PWMdut_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i0.GSR = "DISABLED";
    LUT4 i3095_3_lut (.A(n3844), .B(n1065), .C(addOut[19]), .Z(intgOut0_28__N_1627[19])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3095_3_lut.init = 16'h3232;
    LUT4 mux_1198_i2_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[1]), 
         .D(speed_set_m3[1]), .Z(n5322)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i19_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[18]), 
         .D(speed_set_m3[18]), .Z(n5356)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i16_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[15]), 
         .D(speed_set_m3[15]), .Z(n5350)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i15_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[14]), 
         .D(speed_set_m3[14]), .Z(n5348)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3093_3_lut (.A(n3844), .B(n1065), .C(addOut[16]), .Z(intgOut0_28__N_1627[16])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3093_3_lut.init = 16'h3232;
    LUT4 i3091_3_lut (.A(n3844), .B(n1065), .C(addOut[12]), .Z(intgOut0_28__N_1627[12])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3091_3_lut.init = 16'h3232;
    LUT4 mux_1198_i12_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[11]), 
         .D(speed_set_m3[11]), .Z(n5342)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i20_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[19]), 
         .D(speed_set_m3[19]), .Z(n5358)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17456_4_lut_4_lut_then_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), 
         .D(n22440), .Z(n21731)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 185[26])
    defparam i17456_4_lut_4_lut_then_4_lut.init = 16'hfff7;
    LUT4 mux_1198_i13_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[12]), 
         .D(speed_set_m3[12]), .Z(n5344)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3089_3_lut (.A(n3844), .B(n1065), .C(addOut[11]), .Z(intgOut0_28__N_1627[11])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3089_3_lut.init = 16'h3232;
    LUT4 mux_136_i5_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[4]), 
         .D(backOut1[4]), .Z(n585[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i10_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[9]), 
         .D(backOut1[9]), .Z(n585[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1198_i8_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[7]), 
         .D(speed_set_m3[7]), .Z(n5334)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1198_i6_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[5]), 
         .D(speed_set_m3[5]), .Z(n5330)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_136_i9_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[8]), 
         .D(backOut1[8]), .Z(n585[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1198_i10_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[9]), 
         .D(speed_set_m3[9]), .Z(n5338)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_136_i3_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[2]), 
         .D(backOut1[2]), .Z(n585[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i2_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[1]), 
         .D(backOut1[1]), .Z(n585[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3087_3_lut (.A(n3844), .B(n1065), .C(addOut[10]), .Z(intgOut0_28__N_1627[10])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3087_3_lut.init = 16'h3232;
    LUT4 mux_136_i13_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[12]), 
         .D(backOut1[12]), .Z(n585[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i12_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[11]), 
         .D(backOut1[11]), .Z(n585[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i11_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[10]), 
         .D(backOut1[10]), .Z(n585[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i8_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[7]), 
         .D(backOut1[7]), .Z(n585[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1198_i21_3_lut_4_lut (.A(n16309), .B(n42), .C(speed_set_m2[20]), 
         .D(speed_set_m3[20]), .Z(n5360)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1198_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_323 (.A(subIn1_24__N_1342), .B(n35), .Z(n21636)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam i1_2_lut_rep_323.init = 16'h8888;
    LUT4 mux_136_i6_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[5]), 
         .D(backOut1[5]), .Z(n585[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i4_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[3]), 
         .D(backOut1[3]), .Z(n585[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i14_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[13]), 
         .D(backOut1[13]), .Z(n585[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i16_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m4[15]), .Z(n5392)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1197_i20_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m4[19]), .Z(n5400)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1197_i4_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m4[3]), .Z(n5368)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i7_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[6]), 
         .D(backOut1[6]), .Z(n585[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3085_3_lut (.A(n3844), .B(n1065), .C(addOut[7]), .Z(intgOut0_28__N_1627[7])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3085_3_lut.init = 16'h3232;
    LUT4 mux_136_i15_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[14]), 
         .D(backOut1[14]), .Z(n585[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13273_2_lut (.A(addOut[19]), .B(n22440), .Z(backOut3_28__N_1872[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13273_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_adj_50 (.A(n22440), .B(ss[1]), .Z(n19967)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_adj_50.init = 16'heeee;
    LUT4 i1_4_lut (.A(n16477), .B(n19913), .C(n21677), .D(n22440), .Z(clk_N_875_enable_392)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;
    defparam i1_4_lut.init = 16'hf5dd;
    LUT4 mux_1197_i3_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m4[2]), .Z(n5366)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i16_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[15]), 
         .D(backOut1[15]), .Z(n585[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i17_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[16]), 
         .D(backOut1[16]), .Z(n585[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i2_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m4[1]), .Z(n5364)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i18_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[17]), 
         .D(backOut1[17]), .Z(n585[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i19_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[18]), 
         .D(backOut1[18]), .Z(n585[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i19_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15369_5 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18778), .COUT(n18779));
    defparam add_15369_5.INIT0 = 16'h0aaa;
    defparam add_15369_5.INIT1 = 16'h0aaa;
    defparam add_15369_5.INJECT1_0 = "NO";
    defparam add_15369_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_51 (.A(n3660), .B(n35_adj_2328), .C(n40), .D(n36), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_51.init = 16'haaa8;
    LUT4 mux_136_i20_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[19]), 
         .D(backOut1[19]), .Z(n585[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i1_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m4[0]), .Z(n5320)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i21_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[20]), 
         .D(backOut1[20]), .Z(n585[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i22_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[21]), 
         .D(backOut1[21]), .Z(n585[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 i14_4_lut (.A(speed_set_m2[13]), .B(speed_set_m2[1]), .C(speed_set_m2[12]), 
         .D(speed_set_m2[2]), .Z(n35_adj_2328)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(speed_set_m2[15]), .B(n38), .C(n32), .D(speed_set_m2[10]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 mux_136_i1_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[0]), 
         .D(backOut1[0]), .Z(n585[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 i15_4_lut (.A(speed_set_m2[0]), .B(speed_set_m2[7]), .C(speed_set_m2[17]), 
         .D(speed_set_m2[11]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(speed_set_m2[8]), .B(n34), .C(n24), .D(speed_set_m2[16]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(speed_set_m2[6]), .B(speed_set_m2[3]), .C(speed_set_m2[14]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(speed_set_m2[20]), .B(speed_set_m2[19]), .C(speed_set_m2[9]), 
         .D(speed_set_m2[4]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(speed_set_m2[18]), .B(speed_set_m2[5]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 mux_1197_i19_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m4[18]), .Z(n5398)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i23_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[22]), 
         .D(backOut1[22]), .Z(n585[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i24_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[23]), 
         .D(backOut1[23]), .Z(n585[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i21_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m4[20]), .Z(n5402)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i25_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[24]), 
         .D(backOut1[24]), .Z(n585[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i26_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[25]), 
         .D(backOut1[25]), .Z(n585[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i27_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[26]), 
         .D(backOut1[26]), .Z(n585[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i18_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m4[17]), .Z(n5396)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_92_i13_3_lut (.A(\speed_avg_m3[12] ), .B(\speed_avg_m2[12] ), 
         .C(n22423), .Z(subIn2_24__N_1534[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i13_3_lut.init = 16'hcaca;
    LUT4 mux_136_i28_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[27]), 
         .D(backOut1[27]), .Z(n585[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i29_3_lut_4_lut (.A(n21721), .B(n21684), .C(backOut0[28]), 
         .D(backOut1[28]), .Z(n585[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11647_3_lut_4_lut (.A(n21678), .B(n21628), .C(ss[1]), .D(clk_N_875_enable_389), 
         .Z(n14232)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11647_3_lut_4_lut.init = 16'hfe00;
    LUT4 mux_1197_i13_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m4[12]), .Z(n5386)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i11675_3_lut_4_lut (.A(n21678), .B(n21628), .C(ss[1]), .D(clk_N_875_enable_392), 
         .Z(n14260)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11675_3_lut_4_lut.init = 16'hef00;
    LUT4 mux_139_i13_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[12]), 
         .D(n645[12]), .Z(n675[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i17_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[16]), 
         .D(n645[16]), .Z(n675[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i14_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[13]), 
         .D(n645[13]), .Z(n675[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_adj_52 (.A(n1357[15]), .B(n2297[3]), .C(n30_adj_2327), 
         .Z(n1539[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_52.init = 16'h8a8a;
    LUT4 mux_139_i25_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[24]), 
         .D(n645[24]), .Z(n675[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i6_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m4[5]), .Z(n5372)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1197_i10_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m4[9]), .Z(n5380)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1197_i15_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m4[14]), .Z(n5390)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1197_i12_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m4[11]), .Z(n5384)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_139_i23_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[22]), 
         .D(n645[22]), .Z(n675[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i10_3_lut (.A(\speed_avg_m3[9] ), .B(\speed_avg_m2[9] ), 
         .C(n22423), .Z(subIn2_24__N_1534[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i10_3_lut.init = 16'hcaca;
    LUT4 mux_139_i20_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[19]), 
         .D(n645[19]), .Z(n675[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i12_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[11]), 
         .D(n645[11]), .Z(n675[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i10_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[9]), 
         .D(n645[9]), .Z(n675[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17456_4_lut_4_lut_else_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), 
         .D(n22440), .Z(n21730)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 185[26])
    defparam i17456_4_lut_4_lut_else_4_lut.init = 16'hffb7;
    LUT4 mux_92_i9_3_lut (.A(\speed_avg_m3[8] ), .B(\speed_avg_m2[8] ), 
         .C(n22423), .Z(subIn2_24__N_1534[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i9_3_lut.init = 16'hcaca;
    LUT4 mux_139_i6_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[5]), 
         .D(n645[5]), .Z(n675[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i8_3_lut (.A(\speed_avg_m3[7] ), .B(\speed_avg_m2[7] ), 
         .C(n22423), .Z(subIn2_24__N_1534[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i8_3_lut.init = 16'hcaca;
    LUT4 mux_139_i28_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[27]), 
         .D(n645[27]), .Z(n675[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i4_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[3]), 
         .D(n645[3]), .Z(n675[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i3_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[2]), 
         .D(n645[2]), .Z(n675[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i4_3_lut (.A(\speed_avg_m3[3] ), .B(\speed_avg_m2[3] ), 
         .C(n22423), .Z(subIn2_24__N_1534[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i4_3_lut.init = 16'hcaca;
    LUT4 mux_92_i20_4_lut (.A(\speed_avg_m4[19] ), .B(\speed_avg_m3[19] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i20_4_lut.init = 16'hcac0;
    LUT4 mux_139_i2_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[1]), 
         .D(n645[1]), .Z(n675[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i21_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[20]), 
         .D(n645[20]), .Z(n675[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i18_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[17]), 
         .D(n645[17]), .Z(n675[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i19_4_lut (.A(\speed_avg_m4[18] ), .B(\speed_avg_m3[18] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i19_4_lut.init = 16'hcac0;
    LUT4 mux_139_i16_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[15]), 
         .D(n645[15]), .Z(n675[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i11_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m4[10]), .Z(n5382)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_92_i18_4_lut (.A(\speed_avg_m4[17] ), .B(\speed_avg_m3[17] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i18_4_lut.init = 16'hcac0;
    LUT4 mux_1197_i8_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m4[7]), .Z(n5376)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i13_4_lut_adj_53 (.A(speed_set_m3[20]), .B(speed_set_m3[19]), .C(speed_set_m3[9]), 
         .D(speed_set_m3[4]), .Z(n34_adj_2329)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_53.init = 16'hfffe;
    LUT4 i13135_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[0]), 
         .D(ss[1]), .Z(intgOut3_28__N_1058[0])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13135_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 mux_92_i17_4_lut (.A(\speed_avg_m4[16] ), .B(\speed_avg_m3[16] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i17_4_lut.init = 16'hcac0;
    LUT4 mux_92_i16_4_lut (.A(\speed_avg_m4[15] ), .B(\speed_avg_m3[15] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i16_4_lut.init = 16'hcac0;
    CCU2D add_1188_11 (.A0(n5428), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5430), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18414), 
          .COUT(n18415), .S0(n2353[9]), .S1(n2353[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_11.INIT0 = 16'hf555;
    defparam add_1188_11.INIT1 = 16'hf555;
    defparam add_1188_11.INJECT1_0 = "NO";
    defparam add_1188_11.INJECT1_1 = "NO";
    CCU2D add_1188_9 (.A0(n5424), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5426), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18413), 
          .COUT(n18414), .S0(n2353[7]), .S1(n2353[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_9.INIT0 = 16'hf555;
    defparam add_1188_9.INIT1 = 16'hf555;
    defparam add_1188_9.INJECT1_0 = "NO";
    defparam add_1188_9.INJECT1_1 = "NO";
    LUT4 mux_92_i15_4_lut (.A(\speed_avg_m4[14] ), .B(\speed_avg_m3[14] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i15_4_lut.init = 16'hcac0;
    CCU2D add_1188_7 (.A0(n5420), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5422), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18412), 
          .COUT(n18413), .S0(n2353[5]), .S1(n2353[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_7.INIT0 = 16'hf555;
    defparam add_1188_7.INIT1 = 16'hf555;
    defparam add_1188_7.INJECT1_0 = "NO";
    defparam add_1188_7.INJECT1_1 = "NO";
    LUT4 mux_92_i14_4_lut (.A(\speed_avg_m4[13] ), .B(\speed_avg_m3[13] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i14_4_lut.init = 16'hcac0;
    CCU2D add_1188_5 (.A0(n5416), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5418), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18411), 
          .COUT(n18412), .S0(n2353[3]), .S1(n2353[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_5.INIT0 = 16'hf555;
    defparam add_1188_5.INIT1 = 16'hf555;
    defparam add_1188_5.INJECT1_0 = "NO";
    defparam add_1188_5.INJECT1_1 = "NO";
    CCU2D add_1188_3 (.A0(n5412), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5414), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18410), 
          .COUT(n18411), .S0(n2353[1]), .S1(n2353[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_3.INIT0 = 16'hf555;
    defparam add_1188_3.INIT1 = 16'hf555;
    defparam add_1188_3.INJECT1_0 = "NO";
    defparam add_1188_3.INJECT1_1 = "NO";
    CCU2D add_1182_5 (.A0(n1294[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1294[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18406), 
          .COUT(n18407), .S0(n2261[3]), .S1(n2261[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1182_5.INIT0 = 16'hf555;
    defparam add_1182_5.INIT1 = 16'hf555;
    defparam add_1182_5.INJECT1_0 = "NO";
    defparam add_1182_5.INJECT1_1 = "NO";
    LUT4 mux_92_i12_4_lut (.A(\speed_avg_m4[11] ), .B(\speed_avg_m3[11] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i12_4_lut.init = 16'hcac0;
    LUT4 mux_92_i11_4_lut (.A(\speed_avg_m4[10] ), .B(\speed_avg_m3[10] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i11_4_lut.init = 16'hcac0;
    CCU2D add_1182_9 (.A0(n1294[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1294[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18408), 
          .COUT(n18409), .S0(n2261[7]), .S1(n2261[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1182_9.INIT0 = 16'hf555;
    defparam add_1182_9.INIT1 = 16'hf555;
    defparam add_1182_9.INJECT1_0 = "NO";
    defparam add_1182_9.INJECT1_1 = "NO";
    CCU2D add_1182_3 (.A0(n1294[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1294[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18405), 
          .COUT(n18406), .S0(n2261[1]), .S1(n2261[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1182_3.INIT0 = 16'hf555;
    defparam add_1182_3.INIT1 = 16'hf555;
    defparam add_1182_3.INJECT1_0 = "NO";
    defparam add_1182_3.INJECT1_1 = "NO";
    CCU2D add_1188_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5410), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18410), 
          .S1(n2353[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_1.INIT0 = 16'hF000;
    defparam add_1188_1.INIT1 = 16'h0aaa;
    defparam add_1188_1.INJECT1_0 = "NO";
    defparam add_1188_1.INJECT1_1 = "NO";
    CCU2D add_1182_7 (.A0(n1294[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1294[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18407), 
          .COUT(n18408), .S0(n2261[5]), .S1(n2261[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1182_7.INIT0 = 16'hf555;
    defparam add_1182_7.INIT1 = 16'hf555;
    defparam add_1182_7.INJECT1_0 = "NO";
    defparam add_1182_7.INJECT1_1 = "NO";
    LUT4 i3_2_lut_adj_54 (.A(speed_set_m3[18]), .B(speed_set_m3[5]), .Z(n24_adj_2330)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_54.init = 16'heeee;
    CCU2D add_1182_11 (.A0(n1294[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18409), 
          .S0(n2261[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1182_11.INIT0 = 16'hf555;
    defparam add_1182_11.INIT1 = 16'h0000;
    defparam add_1182_11.INJECT1_0 = "NO";
    defparam add_1182_11.INJECT1_1 = "NO";
    CCU2D add_1182_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1294[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18405), 
          .S1(n2261[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1182_1.INIT0 = 16'hF000;
    defparam add_1182_1.INIT1 = 16'h0aaa;
    defparam add_1182_1.INJECT1_0 = "NO";
    defparam add_1182_1.INJECT1_1 = "NO";
    LUT4 mux_1197_i7_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m4[6]), .Z(n5374)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_92_i7_4_lut (.A(\speed_avg_m4[6] ), .B(\speed_avg_m3[6] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i7_4_lut.init = 16'hcac0;
    LUT4 mux_139_i7_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[6]), 
         .D(n645[6]), .Z(n675[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i7_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX dirout_m2_347 (.D(subIn1_24__N_1533), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m2_347.GSR = "DISABLED";
    FD1P3AX dirout_m3_348 (.D(dirout_m3_N_1947), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m3_348.GSR = "DISABLED";
    FD1P3AX dirout_m1_346 (.D(subIn1_24__N_1347), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m1_346.GSR = "DISABLED";
    FD1P3AX dirout_m4_349 (.D(dirout_m4_N_1950), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m4_349.GSR = "DISABLED";
    LUT4 mux_92_i6_4_lut (.A(\speed_avg_m4[5] ), .B(\speed_avg_m3[5] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i6_4_lut.init = 16'hcac0;
    FD1P3AX backOut1_i0_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i28.GSR = "DISABLED";
    LUT4 mux_92_i5_4_lut (.A(\speed_avg_m4[4] ), .B(\speed_avg_m3[4] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i5_4_lut.init = 16'hcac0;
    CCU2D add_15369_3 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18777), .COUT(n18778));
    defparam add_15369_3.INIT0 = 16'hf555;
    defparam add_15369_3.INIT1 = 16'hf555;
    defparam add_15369_3.INJECT1_0 = "NO";
    defparam add_15369_3.INJECT1_1 = "NO";
    CCU2D add_15369_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[4]), .B1(speed_set_m4[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18777));
    defparam add_15369_1.INIT0 = 16'hF000;
    defparam add_15369_1.INIT1 = 16'ha666;
    defparam add_15369_1.INJECT1_0 = "NO";
    defparam add_15369_1.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_5 (.A0(n2353[3]), .B0(n4425), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[4]), .B1(n4424), .C1(GND_net), .D1(GND_net), 
          .CIN(n18658), .COUT(n18659), .S0(n4472), .S1(n4471));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_5.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_5.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_5.INJECT1_1 = "NO";
    LUT4 mux_92_i3_4_lut (.A(\speed_avg_m4[2] ), .B(\speed_avg_m3[2] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i3_4_lut.init = 16'hcac0;
    FD1P3AX backOut1_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i24.GSR = "DISABLED";
    LUT4 mux_92_i2_4_lut (.A(\speed_avg_m4[1] ), .B(\speed_avg_m3[1] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i2_4_lut.init = 16'hcac0;
    LUT4 mux_92_i1_4_lut (.A(\speed_avg_m4[0] ), .B(\speed_avg_m3[0] ), 
         .C(n21668), .D(n4358), .Z(subIn2_24__N_1534[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i1_4_lut.init = 16'hcac0;
    FD1P3AX backOut1_i0_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i20.GSR = "DISABLED";
    LUT4 mux_1197_i5_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m4[4]), .Z(n5370)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_135_i9_4_lut (.A(backOut2[8]), .B(backOut3[8]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i9_4_lut.init = 16'h0aca;
    FD1P3AX backOut1_i0_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i18.GSR = "DISABLED";
    LUT4 mux_1197_i17_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m4[16]), .Z(n5394)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i17_3_lut_4_lut.init = 16'hf780;
    FD1P3AX backOut1_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i11.GSR = "DISABLED";
    LUT4 mux_139_i24_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[23]), 
         .D(n645[23]), .Z(n675[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i24_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX backOut1_i0_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_44), 
            .CK(clk_N_875), .Q(backOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i1.GSR = "DISABLED";
    LUT4 mux_139_i22_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[21]), 
         .D(n645[21]), .Z(n675[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i19_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[18]), 
         .D(n645[18]), .Z(n675[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13242_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[1]), 
         .D(ss[1]), .Z(intgOut3_28__N_1058[1])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13242_2_lut_3_lut_4_lut.init = 16'h1000;
    CCU2D add_223_13 (.A0(Out3[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18450), 
          .COUT(n18451), .S0(n1357[11]), .S1(n1357[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_13.INIT0 = 16'h5aaa;
    defparam add_223_13.INIT1 = 16'h5aaa;
    defparam add_223_13.INJECT1_0 = "NO";
    defparam add_223_13.INJECT1_1 = "NO";
    LUT4 mux_1197_i9_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m4[8]), .Z(n5378)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_135_i10_4_lut (.A(backOut2[9]), .B(backOut3[9]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i10_4_lut.init = 16'h0aca;
    LUT4 mux_139_i5_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[4]), 
         .D(n645[4]), .Z(n675[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i11_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[10]), 
         .D(n645[10]), .Z(n675[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i29_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[28]), 
         .D(n645[28]), .Z(n675[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i9_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[8]), 
         .D(n645[8]), .Z(n675[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i15_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[14]), 
         .D(n645[14]), .Z(n675[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1197_i14_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m4[13]), .Z(n5388)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1197_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 ss_4__I_0_358_i6_2_lut (.A(ss[0]), .B(ss[1]), .Z(n6)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam ss_4__I_0_358_i6_2_lut.init = 16'hdddd;
    LUT4 mux_139_i26_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[25]), 
         .D(n645[25]), .Z(n675[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_55 (.A(n16473), .B(n19945), .C(n21677), .D(n22440), 
         .Z(clk_N_875_enable_309)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;
    defparam i1_4_lut_adj_55.init = 16'hf5dd;
    LUT4 i13744_2_lut_rep_324 (.A(n16309), .B(n42), .Z(n21637)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13744_2_lut_rep_324.init = 16'heeee;
    LUT4 i13243_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[2]), 
         .D(ss[1]), .Z(intgOut3_28__N_1058[2])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13243_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 mux_135_i11_4_lut (.A(backOut2[10]), .B(backOut3[10]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i11_4_lut.init = 16'h0aca;
    LUT4 mux_139_i27_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[26]), 
         .D(n645[26]), .Z(n675[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i8_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[7]), 
         .D(n645[7]), .Z(n675[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i1_3_lut_4_lut (.A(n21721), .B(n21686), .C(intgOut0[0]), 
         .D(n645[0]), .Z(n675[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13893_3_lut_4_lut (.A(n6), .B(n21686), .C(n4_adj_2332), .D(n3780), 
         .Z(n16473)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13893_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_4_lut_adj_56 (.A(n3756), .B(n35_adj_2333), .C(n40_adj_2334), 
         .D(n36_adj_2335), .Z(n4_adj_2332)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_56.init = 16'haaa8;
    LUT4 i14_4_lut_adj_57 (.A(speed_set_m4[13]), .B(speed_set_m4[1]), .C(speed_set_m4[12]), 
         .D(speed_set_m4[2]), .Z(n35_adj_2333)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_57.init = 16'hfffe;
    LUT4 i19_4_lut_adj_58 (.A(speed_set_m4[15]), .B(n38_adj_2336), .C(n32_adj_2337), 
         .D(speed_set_m4[10]), .Z(n40_adj_2334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_58.init = 16'hfffe;
    LUT4 i15_4_lut_adj_59 (.A(speed_set_m4[0]), .B(speed_set_m4[7]), .C(speed_set_m4[17]), 
         .D(speed_set_m4[11]), .Z(n36_adj_2335)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_59.init = 16'hfffe;
    LUT4 i13889_3_lut_4_lut (.A(n6), .B(n21686), .C(n4_adj_2338), .D(n3732), 
         .Z(n16469)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13889_3_lut_4_lut.init = 16'hfeee;
    LUT4 i17_4_lut_adj_60 (.A(speed_set_m4[8]), .B(n34_adj_2339), .C(n24_adj_2340), 
         .D(speed_set_m4[16]), .Z(n38_adj_2336)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_60.init = 16'hfffe;
    LUT4 mux_135_i12_4_lut (.A(backOut2[11]), .B(backOut3[11]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i12_4_lut.init = 16'h0aca;
    FD1S3AX addOut_2102__i0 (.D(n121[0]), .CK(clk_N_875), .Q(addOut[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i0.GSR = "ENABLED";
    AND2 AND2_t64 (.A(subOut[0]), .B(n21660), .Z(multOut_28__N_1411[0])) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1256[10:66])
    AND2 AND2_t61 (.A(subOut[0]), .B(multIn2[2]), .Z(mult_29s_25s_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1262[10:66])
    AND2 AND2_t58 (.A(subOut[0]), .B(multIn2[8]), .Z(mult_29s_25s_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1268[10:66])
    AND2 AND2_t55 (.A(subOut[0]), .B(multIn2[8]), .Z(mult_29s_25s_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1274[10:66])
    AND2 AND2_t52 (.A(subOut[0]), .B(multIn2[8]), .Z(mult_29s_25s_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1280[10:66])
    AND2 AND2_t49 (.A(subOut[0]), .B(multIn2[10]), .Z(mult_29s_25s_0_pp_5_10)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1286[10:68])
    AND2 AND2_t46 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_6_12)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1292[10:68])
    AND2 AND2_t43 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_7_14)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1298[10:68])
    AND2 AND2_t40 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_8_16)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1304[10:68])
    AND2 AND2_t37 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_9_18)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1310[10:68])
    AND2 AND2_t34 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_10_20)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1316[10:69])
    AND2 AND2_t31 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_11_22)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1322[10:69])
    ND2 ND2_t28 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t27 (.A(subOut[1]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_25)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t26 (.A(subOut[2]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t25 (.A(subOut[3]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_27)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t24 (.A(subOut[4]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i11_3_lut_adj_61 (.A(speed_set_m4[6]), .B(speed_set_m4[3]), .C(speed_set_m4[14]), 
         .Z(n32_adj_2337)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_61.init = 16'hfefe;
    FADD2B mult_29s_25s_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_12 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_14 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_16 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_18 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_20 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_22 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_0_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_0_2), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_1_2), .CI(GND_net), .COUT(co_mult_29s_25s_0_0_1), 
           .S1(multOut_28__N_1411[2])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_2 (.A0(mult_29s_25s_0_pp_0_3), .A1(mult_29s_25s_0_pp_0_4), 
           .B0(mult_29s_25s_0_pp_1_3), .B1(mult_29s_25s_0_pp_1_4), .CI(co_mult_29s_25s_0_0_1), 
           .COUT(co_mult_29s_25s_0_0_2), .S0(multOut_28__N_1411[3]), .S1(s_mult_29s_25s_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_3 (.A0(mult_29s_25s_0_pp_0_5), .A1(mult_29s_25s_0_pp_0_6), 
           .B0(mult_29s_25s_0_pp_1_5), .B1(mult_29s_25s_0_pp_1_6), .CI(co_mult_29s_25s_0_0_2), 
           .COUT(co_mult_29s_25s_0_0_3), .S0(s_mult_29s_25s_0_0_5), .S1(s_mult_29s_25s_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_4 (.A0(mult_29s_25s_0_pp_0_7), .A1(mult_29s_25s_0_pp_0_8), 
           .B0(mult_29s_25s_0_pp_1_7), .B1(mult_29s_25s_0_pp_1_8), .CI(co_mult_29s_25s_0_0_3), 
           .COUT(co_mult_29s_25s_0_0_4), .S0(s_mult_29s_25s_0_0_7), .S1(s_mult_29s_25s_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_5 (.A0(mult_29s_25s_0_pp_0_9), .A1(mult_29s_25s_0_pp_0_10), 
           .B0(mult_29s_25s_0_pp_1_9), .B1(mult_29s_25s_0_pp_1_10), .CI(co_mult_29s_25s_0_0_4), 
           .COUT(co_mult_29s_25s_0_0_5), .S0(s_mult_29s_25s_0_0_9), .S1(s_mult_29s_25s_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_6 (.A0(mult_29s_25s_0_pp_0_11), .A1(mult_29s_25s_0_pp_0_12), 
           .B0(mult_29s_25s_0_pp_1_11), .B1(mult_29s_25s_0_pp_1_12), .CI(co_mult_29s_25s_0_0_5), 
           .COUT(co_mult_29s_25s_0_0_6), .S0(s_mult_29s_25s_0_0_11), .S1(s_mult_29s_25s_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_7 (.A0(mult_29s_25s_0_pp_0_13), .A1(mult_29s_25s_0_pp_0_14), 
           .B0(mult_29s_25s_0_pp_1_13), .B1(mult_29s_25s_0_pp_1_14), .CI(co_mult_29s_25s_0_0_6), 
           .COUT(co_mult_29s_25s_0_0_7), .S0(s_mult_29s_25s_0_0_13), .S1(s_mult_29s_25s_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_8 (.A0(mult_29s_25s_0_pp_0_15), .A1(mult_29s_25s_0_pp_0_16), 
           .B0(mult_29s_25s_0_pp_1_15), .B1(mult_29s_25s_0_pp_1_16), .CI(co_mult_29s_25s_0_0_7), 
           .COUT(co_mult_29s_25s_0_0_8), .S0(s_mult_29s_25s_0_0_15), .S1(s_mult_29s_25s_0_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_9 (.A0(mult_29s_25s_0_pp_0_17), .A1(mult_29s_25s_0_pp_0_18), 
           .B0(mult_29s_25s_0_pp_1_17), .B1(mult_29s_25s_0_pp_1_18), .CI(co_mult_29s_25s_0_0_8), 
           .COUT(co_mult_29s_25s_0_0_9), .S0(s_mult_29s_25s_0_0_17), .S1(s_mult_29s_25s_0_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_10 (.A0(mult_29s_25s_0_pp_0_19), .A1(mult_29s_25s_0_pp_0_20), 
           .B0(mult_29s_25s_0_pp_1_19), .B1(mult_29s_25s_0_pp_1_20), .CI(co_mult_29s_25s_0_0_9), 
           .COUT(co_mult_29s_25s_0_0_10), .S0(s_mult_29s_25s_0_0_19), .S1(s_mult_29s_25s_0_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_11 (.A0(mult_29s_25s_0_pp_0_21), .A1(mult_29s_25s_0_pp_0_22), 
           .B0(mult_29s_25s_0_pp_1_21), .B1(mult_29s_25s_0_pp_1_22), .CI(co_mult_29s_25s_0_0_10), 
           .COUT(co_mult_29s_25s_0_0_11), .S0(s_mult_29s_25s_0_0_21), .S1(s_mult_29s_25s_0_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_12 (.A0(mult_29s_25s_0_pp_0_23), .A1(mult_29s_25s_0_pp_0_24), 
           .B0(mult_29s_25s_0_pp_1_23), .B1(mult_29s_25s_0_pp_1_24), .CI(co_mult_29s_25s_0_0_11), 
           .COUT(co_mult_29s_25s_0_0_12), .S0(s_mult_29s_25s_0_0_23), .S1(s_mult_29s_25s_0_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_13 (.A0(mult_29s_25s_0_pp_0_25), .A1(mult_29s_25s_0_pp_0_26), 
           .B0(mult_29s_25s_0_pp_1_25), .B1(mult_29s_25s_0_pp_1_26), .CI(co_mult_29s_25s_0_0_12), 
           .COUT(co_mult_29s_25s_0_0_13), .S0(s_mult_29s_25s_0_0_25), .S1(s_mult_29s_25s_0_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_14 (.A0(mult_29s_25s_0_pp_0_27), .A1(mult_29s_25s_0_pp_0_28), 
           .B0(mult_29s_25s_0_pp_1_27), .B1(mult_29s_25s_0_pp_1_28), .CI(co_mult_29s_25s_0_0_13), 
           .S0(s_mult_29s_25s_0_0_27), .S1(s_mult_29s_25s_0_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i13901_3_lut_4_lut (.A(n6), .B(n21686), .C(n4_adj_2341), .D(n3636), 
         .Z(n16481)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13901_3_lut_4_lut.init = 16'hfeee;
    FADD2B Cadd_mult_29s_25s_0_1_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_2_6), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_3_6), .CI(GND_net), .COUT(co_mult_29s_25s_0_1_1), 
           .S1(s_mult_29s_25s_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_2 (.A0(mult_29s_25s_0_pp_2_7), .A1(mult_29s_25s_0_pp_2_8), 
           .B0(mult_29s_25s_0_pp_3_7), .B1(mult_29s_25s_0_pp_3_8), .CI(co_mult_29s_25s_0_1_1), 
           .COUT(co_mult_29s_25s_0_1_2), .S0(s_mult_29s_25s_0_1_7), .S1(s_mult_29s_25s_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_3 (.A0(mult_29s_25s_0_pp_2_9), .A1(mult_29s_25s_0_pp_2_10), 
           .B0(mult_29s_25s_0_pp_3_9), .B1(mult_29s_25s_0_pp_3_10), .CI(co_mult_29s_25s_0_1_2), 
           .COUT(co_mult_29s_25s_0_1_3), .S0(s_mult_29s_25s_0_1_9), .S1(s_mult_29s_25s_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_4 (.A0(mult_29s_25s_0_pp_2_11), .A1(mult_29s_25s_0_pp_2_12), 
           .B0(mult_29s_25s_0_pp_3_11), .B1(mult_29s_25s_0_pp_3_12), .CI(co_mult_29s_25s_0_1_3), 
           .COUT(co_mult_29s_25s_0_1_4), .S0(s_mult_29s_25s_0_1_11), .S1(s_mult_29s_25s_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_5 (.A0(mult_29s_25s_0_pp_2_13), .A1(mult_29s_25s_0_pp_2_14), 
           .B0(mult_29s_25s_0_pp_3_13), .B1(mult_29s_25s_0_pp_3_14), .CI(co_mult_29s_25s_0_1_4), 
           .COUT(co_mult_29s_25s_0_1_5), .S0(s_mult_29s_25s_0_1_13), .S1(s_mult_29s_25s_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_6 (.A0(mult_29s_25s_0_pp_2_15), .A1(mult_29s_25s_0_pp_2_16), 
           .B0(mult_29s_25s_0_pp_3_15), .B1(mult_29s_25s_0_pp_3_16), .CI(co_mult_29s_25s_0_1_5), 
           .COUT(co_mult_29s_25s_0_1_6), .S0(s_mult_29s_25s_0_1_15), .S1(s_mult_29s_25s_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_7 (.A0(mult_29s_25s_0_pp_2_17), .A1(mult_29s_25s_0_pp_2_18), 
           .B0(mult_29s_25s_0_pp_3_17), .B1(mult_29s_25s_0_pp_3_18), .CI(co_mult_29s_25s_0_1_6), 
           .COUT(co_mult_29s_25s_0_1_7), .S0(s_mult_29s_25s_0_1_17), .S1(s_mult_29s_25s_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_8 (.A0(mult_29s_25s_0_pp_2_19), .A1(mult_29s_25s_0_pp_2_20), 
           .B0(mult_29s_25s_0_pp_3_19), .B1(mult_29s_25s_0_pp_3_20), .CI(co_mult_29s_25s_0_1_7), 
           .COUT(co_mult_29s_25s_0_1_8), .S0(s_mult_29s_25s_0_1_19), .S1(s_mult_29s_25s_0_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_9 (.A0(mult_29s_25s_0_pp_2_21), .A1(mult_29s_25s_0_pp_2_22), 
           .B0(mult_29s_25s_0_pp_3_21), .B1(mult_29s_25s_0_pp_3_22), .CI(co_mult_29s_25s_0_1_8), 
           .COUT(co_mult_29s_25s_0_1_9), .S0(s_mult_29s_25s_0_1_21), .S1(s_mult_29s_25s_0_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_10 (.A0(mult_29s_25s_0_pp_2_23), .A1(mult_29s_25s_0_pp_2_24), 
           .B0(mult_29s_25s_0_pp_3_23), .B1(mult_29s_25s_0_pp_3_24), .CI(co_mult_29s_25s_0_1_9), 
           .COUT(co_mult_29s_25s_0_1_10), .S0(s_mult_29s_25s_0_1_23), .S1(s_mult_29s_25s_0_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_11 (.A0(mult_29s_25s_0_pp_2_25), .A1(mult_29s_25s_0_pp_2_26), 
           .B0(mult_29s_25s_0_pp_3_25), .B1(mult_29s_25s_0_pp_3_26), .CI(co_mult_29s_25s_0_1_10), 
           .COUT(co_mult_29s_25s_0_1_11), .S0(s_mult_29s_25s_0_1_25), .S1(s_mult_29s_25s_0_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_12 (.A0(mult_29s_25s_0_pp_2_27), .A1(mult_29s_25s_0_pp_2_28), 
           .B0(mult_29s_25s_0_pp_3_27), .B1(mult_29s_25s_0_pp_3_28), .CI(co_mult_29s_25s_0_1_11), 
           .S0(s_mult_29s_25s_0_1_27), .S1(s_mult_29s_25s_0_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_2_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_4_10), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_5_10), .CI(GND_net), .COUT(co_mult_29s_25s_0_2_1), 
           .S1(s_mult_29s_25s_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_2 (.A0(mult_29s_25s_0_pp_4_11), .A1(mult_29s_25s_0_pp_4_12), 
           .B0(mult_29s_25s_0_pp_5_11), .B1(mult_29s_25s_0_pp_5_12), .CI(co_mult_29s_25s_0_2_1), 
           .COUT(co_mult_29s_25s_0_2_2), .S0(s_mult_29s_25s_0_2_11), .S1(s_mult_29s_25s_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_3 (.A0(mult_29s_25s_0_pp_4_13), .A1(mult_29s_25s_0_pp_4_14), 
           .B0(mult_29s_25s_0_pp_5_13), .B1(mult_29s_25s_0_pp_5_14), .CI(co_mult_29s_25s_0_2_2), 
           .COUT(co_mult_29s_25s_0_2_3), .S0(s_mult_29s_25s_0_2_13), .S1(s_mult_29s_25s_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_4 (.A0(mult_29s_25s_0_pp_4_15), .A1(mult_29s_25s_0_pp_4_16), 
           .B0(mult_29s_25s_0_pp_5_15), .B1(mult_29s_25s_0_pp_5_16), .CI(co_mult_29s_25s_0_2_3), 
           .COUT(co_mult_29s_25s_0_2_4), .S0(s_mult_29s_25s_0_2_15), .S1(s_mult_29s_25s_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_5 (.A0(mult_29s_25s_0_pp_4_17), .A1(mult_29s_25s_0_pp_4_18), 
           .B0(mult_29s_25s_0_pp_5_17), .B1(mult_29s_25s_0_pp_5_18), .CI(co_mult_29s_25s_0_2_4), 
           .COUT(co_mult_29s_25s_0_2_5), .S0(s_mult_29s_25s_0_2_17), .S1(s_mult_29s_25s_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_6 (.A0(mult_29s_25s_0_pp_4_19), .A1(mult_29s_25s_0_pp_4_20), 
           .B0(mult_29s_25s_0_pp_5_19), .B1(mult_29s_25s_0_pp_5_20), .CI(co_mult_29s_25s_0_2_5), 
           .COUT(co_mult_29s_25s_0_2_6), .S0(s_mult_29s_25s_0_2_19), .S1(s_mult_29s_25s_0_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_7 (.A0(mult_29s_25s_0_pp_4_21), .A1(mult_29s_25s_0_pp_4_22), 
           .B0(mult_29s_25s_0_pp_5_21), .B1(mult_29s_25s_0_pp_5_22), .CI(co_mult_29s_25s_0_2_6), 
           .COUT(co_mult_29s_25s_0_2_7), .S0(s_mult_29s_25s_0_2_21), .S1(s_mult_29s_25s_0_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_8 (.A0(mult_29s_25s_0_pp_4_23), .A1(mult_29s_25s_0_pp_4_24), 
           .B0(mult_29s_25s_0_pp_5_23), .B1(mult_29s_25s_0_pp_5_24), .CI(co_mult_29s_25s_0_2_7), 
           .COUT(co_mult_29s_25s_0_2_8), .S0(s_mult_29s_25s_0_2_23), .S1(s_mult_29s_25s_0_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_9 (.A0(mult_29s_25s_0_pp_4_25), .A1(mult_29s_25s_0_pp_4_26), 
           .B0(mult_29s_25s_0_pp_5_25), .B1(mult_29s_25s_0_pp_5_26), .CI(co_mult_29s_25s_0_2_8), 
           .COUT(co_mult_29s_25s_0_2_9), .S0(s_mult_29s_25s_0_2_25), .S1(s_mult_29s_25s_0_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_10 (.A0(mult_29s_25s_0_pp_4_27), .A1(mult_29s_25s_0_pp_4_28), 
           .B0(mult_29s_25s_0_pp_5_27), .B1(mult_29s_25s_0_pp_5_28), .CI(co_mult_29s_25s_0_2_9), 
           .S0(s_mult_29s_25s_0_2_27), .S1(s_mult_29s_25s_0_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i13897_3_lut_4_lut (.A(n6), .B(n21686), .C(n4), .D(n3684), 
         .Z(n16477)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13897_3_lut_4_lut.init = 16'hfeee;
    FADD2B Cadd_mult_29s_25s_0_3_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_6_14), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_7_14), .CI(GND_net), .COUT(co_mult_29s_25s_0_3_1), 
           .S1(s_mult_29s_25s_0_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_2 (.A0(mult_29s_25s_0_pp_6_15), .A1(mult_29s_25s_0_pp_6_16), 
           .B0(mult_29s_25s_0_pp_7_15), .B1(mult_29s_25s_0_pp_7_16), .CI(co_mult_29s_25s_0_3_1), 
           .COUT(co_mult_29s_25s_0_3_2), .S0(s_mult_29s_25s_0_3_15), .S1(s_mult_29s_25s_0_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_3 (.A0(mult_29s_25s_0_pp_6_17), .A1(mult_29s_25s_0_pp_6_18), 
           .B0(mult_29s_25s_0_pp_7_17), .B1(mult_29s_25s_0_pp_7_18), .CI(co_mult_29s_25s_0_3_2), 
           .COUT(co_mult_29s_25s_0_3_3), .S0(s_mult_29s_25s_0_3_17), .S1(s_mult_29s_25s_0_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_4 (.A0(mult_29s_25s_0_pp_6_19), .A1(mult_29s_25s_0_pp_6_20), 
           .B0(mult_29s_25s_0_pp_7_19), .B1(mult_29s_25s_0_pp_7_20), .CI(co_mult_29s_25s_0_3_3), 
           .COUT(co_mult_29s_25s_0_3_4), .S0(s_mult_29s_25s_0_3_19), .S1(s_mult_29s_25s_0_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_5 (.A0(mult_29s_25s_0_pp_6_21), .A1(mult_29s_25s_0_pp_6_22), 
           .B0(mult_29s_25s_0_pp_7_21), .B1(mult_29s_25s_0_pp_7_22), .CI(co_mult_29s_25s_0_3_4), 
           .COUT(co_mult_29s_25s_0_3_5), .S0(s_mult_29s_25s_0_3_21), .S1(s_mult_29s_25s_0_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_6 (.A0(mult_29s_25s_0_pp_6_23), .A1(mult_29s_25s_0_pp_6_24), 
           .B0(mult_29s_25s_0_pp_7_23), .B1(mult_29s_25s_0_pp_7_24), .CI(co_mult_29s_25s_0_3_5), 
           .COUT(co_mult_29s_25s_0_3_6), .S0(s_mult_29s_25s_0_3_23), .S1(s_mult_29s_25s_0_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_7 (.A0(mult_29s_25s_0_pp_6_25), .A1(mult_29s_25s_0_pp_6_26), 
           .B0(mult_29s_25s_0_pp_7_25), .B1(mult_29s_25s_0_pp_7_26), .CI(co_mult_29s_25s_0_3_6), 
           .COUT(co_mult_29s_25s_0_3_7), .S0(s_mult_29s_25s_0_3_25), .S1(s_mult_29s_25s_0_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_8 (.A0(mult_29s_25s_0_pp_6_27), .A1(mult_29s_25s_0_pp_6_28), 
           .B0(mult_29s_25s_0_pp_7_27), .B1(mult_29s_25s_0_pp_7_28), .CI(co_mult_29s_25s_0_3_7), 
           .S0(s_mult_29s_25s_0_3_27), .S1(s_mult_29s_25s_0_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_4_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_8_18), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_9_18), .CI(GND_net), .COUT(co_mult_29s_25s_0_4_1), 
           .S1(s_mult_29s_25s_0_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_2 (.A0(mult_29s_25s_0_pp_8_19), .A1(mult_29s_25s_0_pp_8_20), 
           .B0(mult_29s_25s_0_pp_9_19), .B1(mult_29s_25s_0_pp_9_20), .CI(co_mult_29s_25s_0_4_1), 
           .COUT(co_mult_29s_25s_0_4_2), .S0(s_mult_29s_25s_0_4_19), .S1(s_mult_29s_25s_0_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_3 (.A0(mult_29s_25s_0_pp_8_21), .A1(mult_29s_25s_0_pp_8_22), 
           .B0(mult_29s_25s_0_pp_9_21), .B1(mult_29s_25s_0_pp_9_22), .CI(co_mult_29s_25s_0_4_2), 
           .COUT(co_mult_29s_25s_0_4_3), .S0(s_mult_29s_25s_0_4_21), .S1(s_mult_29s_25s_0_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_4 (.A0(mult_29s_25s_0_pp_8_23), .A1(mult_29s_25s_0_pp_8_24), 
           .B0(mult_29s_25s_0_pp_9_23), .B1(mult_29s_25s_0_pp_9_24), .CI(co_mult_29s_25s_0_4_3), 
           .COUT(co_mult_29s_25s_0_4_4), .S0(s_mult_29s_25s_0_4_23), .S1(s_mult_29s_25s_0_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_5 (.A0(mult_29s_25s_0_pp_8_25), .A1(mult_29s_25s_0_pp_8_26), 
           .B0(mult_29s_25s_0_pp_9_25), .B1(mult_29s_25s_0_pp_9_26), .CI(co_mult_29s_25s_0_4_4), 
           .COUT(co_mult_29s_25s_0_4_5), .S0(s_mult_29s_25s_0_4_25), .S1(s_mult_29s_25s_0_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_6 (.A0(mult_29s_25s_0_pp_8_27), .A1(mult_29s_25s_0_pp_8_28), 
           .B0(mult_29s_25s_0_pp_9_27), .B1(mult_29s_25s_0_pp_9_28), .CI(co_mult_29s_25s_0_4_5), 
           .S0(s_mult_29s_25s_0_4_27), .S1(s_mult_29s_25s_0_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_5_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_10_22), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_11_22), .CI(GND_net), .COUT(co_mult_29s_25s_0_5_1), 
           .S1(s_mult_29s_25s_0_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_2 (.A0(mult_29s_25s_0_pp_10_23), .A1(mult_29s_25s_0_pp_10_24), 
           .B0(mult_29s_25s_0_pp_11_23), .B1(mult_29s_25s_0_pp_11_24), .CI(co_mult_29s_25s_0_5_1), 
           .COUT(co_mult_29s_25s_0_5_2), .S0(s_mult_29s_25s_0_5_23), .S1(s_mult_29s_25s_0_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_3 (.A0(mult_29s_25s_0_pp_10_25), .A1(mult_29s_25s_0_pp_10_26), 
           .B0(mult_29s_25s_0_pp_11_25), .B1(mult_29s_25s_0_pp_11_26), .CI(co_mult_29s_25s_0_5_2), 
           .COUT(co_mult_29s_25s_0_5_3), .S0(s_mult_29s_25s_0_5_25), .S1(s_mult_29s_25s_0_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_4 (.A0(mult_29s_25s_0_pp_10_27), .A1(mult_29s_25s_0_pp_10_28), 
           .B0(mult_29s_25s_0_pp_11_27), .B1(mult_29s_25s_0_pp_11_28), .CI(co_mult_29s_25s_0_5_3), 
           .S0(s_mult_29s_25s_0_5_27), .S1(s_mult_29s_25s_0_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_6_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_12_24), 
           .B0(GND_net), .B1(VCC_net), .CI(GND_net), .COUT(co_mult_29s_25s_0_6_1), 
           .S1(s_mult_29s_25s_0_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_2 (.A0(mult_29s_25s_0_pp_12_25), .A1(mult_29s_25s_0_pp_12_26), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_1), .COUT(co_mult_29s_25s_0_6_2), 
           .S0(s_mult_29s_25s_0_6_25), .S1(s_mult_29s_25s_0_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_3 (.A0(mult_29s_25s_0_pp_12_27), .A1(mult_29s_25s_0_pp_12_28), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_2), .S0(s_mult_29s_25s_0_6_27), 
           .S1(s_mult_29s_25s_0_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i13_4_lut_adj_62 (.A(speed_set_m4[20]), .B(speed_set_m4[19]), .C(speed_set_m4[9]), 
         .D(speed_set_m4[4]), .Z(n34_adj_2339)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_62.init = 16'hfffe;
    FADD2B Cadd_mult_29s_25s_0_7_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_0_4), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_2_4), .CI(GND_net), .COUT(co_mult_29s_25s_0_7_1), 
           .S1(multOut_28__N_1411[4])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_2 (.A0(s_mult_29s_25s_0_0_5), .A1(s_mult_29s_25s_0_0_6), 
           .B0(mult_29s_25s_0_pp_2_5), .B1(s_mult_29s_25s_0_1_6), .CI(co_mult_29s_25s_0_7_1), 
           .COUT(co_mult_29s_25s_0_7_2), .S0(multOut_28__N_1411[5]), .S1(multOut_28__N_1411[6])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_3 (.A0(s_mult_29s_25s_0_0_7), .A1(s_mult_29s_25s_0_0_8), 
           .B0(s_mult_29s_25s_0_1_7), .B1(s_mult_29s_25s_0_1_8), .CI(co_mult_29s_25s_0_7_2), 
           .COUT(co_mult_29s_25s_0_7_3), .S0(multOut_28__N_1411[7]), .S1(s_mult_29s_25s_0_7_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_4 (.A0(s_mult_29s_25s_0_0_9), .A1(s_mult_29s_25s_0_0_10), 
           .B0(s_mult_29s_25s_0_1_9), .B1(s_mult_29s_25s_0_1_10), .CI(co_mult_29s_25s_0_7_3), 
           .COUT(co_mult_29s_25s_0_7_4), .S0(s_mult_29s_25s_0_7_9), .S1(s_mult_29s_25s_0_7_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_5 (.A0(s_mult_29s_25s_0_0_11), .A1(s_mult_29s_25s_0_0_12), 
           .B0(s_mult_29s_25s_0_1_11), .B1(s_mult_29s_25s_0_1_12), .CI(co_mult_29s_25s_0_7_4), 
           .COUT(co_mult_29s_25s_0_7_5), .S0(s_mult_29s_25s_0_7_11), .S1(s_mult_29s_25s_0_7_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_6 (.A0(s_mult_29s_25s_0_0_13), .A1(s_mult_29s_25s_0_0_14), 
           .B0(s_mult_29s_25s_0_1_13), .B1(s_mult_29s_25s_0_1_14), .CI(co_mult_29s_25s_0_7_5), 
           .COUT(co_mult_29s_25s_0_7_6), .S0(s_mult_29s_25s_0_7_13), .S1(s_mult_29s_25s_0_7_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_7 (.A0(s_mult_29s_25s_0_0_15), .A1(s_mult_29s_25s_0_0_16), 
           .B0(s_mult_29s_25s_0_1_15), .B1(s_mult_29s_25s_0_1_16), .CI(co_mult_29s_25s_0_7_6), 
           .COUT(co_mult_29s_25s_0_7_7), .S0(s_mult_29s_25s_0_7_15), .S1(s_mult_29s_25s_0_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_8 (.A0(s_mult_29s_25s_0_0_17), .A1(s_mult_29s_25s_0_0_18), 
           .B0(s_mult_29s_25s_0_1_17), .B1(s_mult_29s_25s_0_1_18), .CI(co_mult_29s_25s_0_7_7), 
           .COUT(co_mult_29s_25s_0_7_8), .S0(s_mult_29s_25s_0_7_17), .S1(s_mult_29s_25s_0_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_9 (.A0(s_mult_29s_25s_0_0_19), .A1(s_mult_29s_25s_0_0_20), 
           .B0(s_mult_29s_25s_0_1_19), .B1(s_mult_29s_25s_0_1_20), .CI(co_mult_29s_25s_0_7_8), 
           .COUT(co_mult_29s_25s_0_7_9), .S0(s_mult_29s_25s_0_7_19), .S1(s_mult_29s_25s_0_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_10 (.A0(s_mult_29s_25s_0_0_21), .A1(s_mult_29s_25s_0_0_22), 
           .B0(s_mult_29s_25s_0_1_21), .B1(s_mult_29s_25s_0_1_22), .CI(co_mult_29s_25s_0_7_9), 
           .COUT(co_mult_29s_25s_0_7_10), .S0(s_mult_29s_25s_0_7_21), .S1(s_mult_29s_25s_0_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_11 (.A0(s_mult_29s_25s_0_0_23), .A1(s_mult_29s_25s_0_0_24), 
           .B0(s_mult_29s_25s_0_1_23), .B1(s_mult_29s_25s_0_1_24), .CI(co_mult_29s_25s_0_7_10), 
           .COUT(co_mult_29s_25s_0_7_11), .S0(s_mult_29s_25s_0_7_23), .S1(s_mult_29s_25s_0_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_12 (.A0(s_mult_29s_25s_0_0_25), .A1(s_mult_29s_25s_0_0_26), 
           .B0(s_mult_29s_25s_0_1_25), .B1(s_mult_29s_25s_0_1_26), .CI(co_mult_29s_25s_0_7_11), 
           .COUT(co_mult_29s_25s_0_7_12), .S0(s_mult_29s_25s_0_7_25), .S1(s_mult_29s_25s_0_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_13 (.A0(s_mult_29s_25s_0_0_27), .A1(s_mult_29s_25s_0_0_28), 
           .B0(s_mult_29s_25s_0_1_27), .B1(s_mult_29s_25s_0_1_28), .CI(co_mult_29s_25s_0_7_12), 
           .S0(s_mult_29s_25s_0_7_27), .S1(s_mult_29s_25s_0_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_8_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_2_12), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_6_12), .CI(GND_net), .COUT(co_mult_29s_25s_0_8_1), 
           .S1(s_mult_29s_25s_0_8_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_2 (.A0(s_mult_29s_25s_0_2_13), .A1(s_mult_29s_25s_0_2_14), 
           .B0(mult_29s_25s_0_pp_6_13), .B1(s_mult_29s_25s_0_3_14), .CI(co_mult_29s_25s_0_8_1), 
           .COUT(co_mult_29s_25s_0_8_2), .S0(s_mult_29s_25s_0_8_13), .S1(s_mult_29s_25s_0_8_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_3 (.A0(s_mult_29s_25s_0_2_15), .A1(s_mult_29s_25s_0_2_16), 
           .B0(s_mult_29s_25s_0_3_15), .B1(s_mult_29s_25s_0_3_16), .CI(co_mult_29s_25s_0_8_2), 
           .COUT(co_mult_29s_25s_0_8_3), .S0(s_mult_29s_25s_0_8_15), .S1(s_mult_29s_25s_0_8_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_4 (.A0(s_mult_29s_25s_0_2_17), .A1(s_mult_29s_25s_0_2_18), 
           .B0(s_mult_29s_25s_0_3_17), .B1(s_mult_29s_25s_0_3_18), .CI(co_mult_29s_25s_0_8_3), 
           .COUT(co_mult_29s_25s_0_8_4), .S0(s_mult_29s_25s_0_8_17), .S1(s_mult_29s_25s_0_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_5 (.A0(s_mult_29s_25s_0_2_19), .A1(s_mult_29s_25s_0_2_20), 
           .B0(s_mult_29s_25s_0_3_19), .B1(s_mult_29s_25s_0_3_20), .CI(co_mult_29s_25s_0_8_4), 
           .COUT(co_mult_29s_25s_0_8_5), .S0(s_mult_29s_25s_0_8_19), .S1(s_mult_29s_25s_0_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_6 (.A0(s_mult_29s_25s_0_2_21), .A1(s_mult_29s_25s_0_2_22), 
           .B0(s_mult_29s_25s_0_3_21), .B1(s_mult_29s_25s_0_3_22), .CI(co_mult_29s_25s_0_8_5), 
           .COUT(co_mult_29s_25s_0_8_6), .S0(s_mult_29s_25s_0_8_21), .S1(s_mult_29s_25s_0_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_7 (.A0(s_mult_29s_25s_0_2_23), .A1(s_mult_29s_25s_0_2_24), 
           .B0(s_mult_29s_25s_0_3_23), .B1(s_mult_29s_25s_0_3_24), .CI(co_mult_29s_25s_0_8_6), 
           .COUT(co_mult_29s_25s_0_8_7), .S0(s_mult_29s_25s_0_8_23), .S1(s_mult_29s_25s_0_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_8 (.A0(s_mult_29s_25s_0_2_25), .A1(s_mult_29s_25s_0_2_26), 
           .B0(s_mult_29s_25s_0_3_25), .B1(s_mult_29s_25s_0_3_26), .CI(co_mult_29s_25s_0_8_7), 
           .COUT(co_mult_29s_25s_0_8_8), .S0(s_mult_29s_25s_0_8_25), .S1(s_mult_29s_25s_0_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_9 (.A0(s_mult_29s_25s_0_2_27), .A1(s_mult_29s_25s_0_2_28), 
           .B0(s_mult_29s_25s_0_3_27), .B1(s_mult_29s_25s_0_3_28), .CI(co_mult_29s_25s_0_8_8), 
           .S0(s_mult_29s_25s_0_8_27), .S1(s_mult_29s_25s_0_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i13759_2_lut_3_lut_4_lut (.A(n16309), .B(n42), .C(n49), .D(n15564), 
         .Z(n16337)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i13759_2_lut_3_lut_4_lut.init = 16'heee0;
    FADD2B Cadd_mult_29s_25s_0_9_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_4_20), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_10_20), .CI(GND_net), .COUT(co_mult_29s_25s_0_9_1), 
           .S1(s_mult_29s_25s_0_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_2 (.A0(s_mult_29s_25s_0_4_21), .A1(s_mult_29s_25s_0_4_22), 
           .B0(mult_29s_25s_0_pp_10_21), .B1(s_mult_29s_25s_0_5_22), .CI(co_mult_29s_25s_0_9_1), 
           .COUT(co_mult_29s_25s_0_9_2), .S0(s_mult_29s_25s_0_9_21), .S1(s_mult_29s_25s_0_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_3 (.A0(s_mult_29s_25s_0_4_23), .A1(s_mult_29s_25s_0_4_24), 
           .B0(s_mult_29s_25s_0_5_23), .B1(s_mult_29s_25s_0_5_24), .CI(co_mult_29s_25s_0_9_2), 
           .COUT(co_mult_29s_25s_0_9_3), .S0(s_mult_29s_25s_0_9_23), .S1(s_mult_29s_25s_0_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_4 (.A0(s_mult_29s_25s_0_4_25), .A1(s_mult_29s_25s_0_4_26), 
           .B0(s_mult_29s_25s_0_5_25), .B1(s_mult_29s_25s_0_5_26), .CI(co_mult_29s_25s_0_9_3), 
           .COUT(co_mult_29s_25s_0_9_4), .S0(s_mult_29s_25s_0_9_25), .S1(s_mult_29s_25s_0_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_5 (.A0(s_mult_29s_25s_0_4_27), .A1(s_mult_29s_25s_0_4_28), 
           .B0(s_mult_29s_25s_0_5_27), .B1(s_mult_29s_25s_0_5_28), .CI(co_mult_29s_25s_0_9_4), 
           .S0(s_mult_29s_25s_0_9_27), .S1(s_mult_29s_25s_0_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i3_2_lut_adj_63 (.A(speed_set_m4[18]), .B(speed_set_m4[5]), .Z(n24_adj_2340)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_63.init = 16'heeee;
    LUT4 subIn2_24__I_25_i13_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[12] ), 
         .D(subIn2_24__N_1534[12]), .Z(subIn2_24__N_1348[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i13_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_mult_29s_25s_0_10_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_7_8), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_4_8), .CI(GND_net), .COUT(co_mult_29s_25s_0_10_1), 
           .S1(multOut_28__N_1411[8])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_2 (.A0(s_mult_29s_25s_0_7_9), .A1(s_mult_29s_25s_0_7_10), 
           .B0(mult_29s_25s_0_pp_4_9), .B1(s_mult_29s_25s_0_2_10), .CI(co_mult_29s_25s_0_10_1), 
           .COUT(co_mult_29s_25s_0_10_2), .S0(multOut_28__N_1411[9]), .S1(multOut_28__N_1411[10])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_3 (.A0(s_mult_29s_25s_0_7_11), .A1(s_mult_29s_25s_0_7_12), 
           .B0(s_mult_29s_25s_0_2_11), .B1(s_mult_29s_25s_0_8_12), .CI(co_mult_29s_25s_0_10_2), 
           .COUT(co_mult_29s_25s_0_10_3), .S0(multOut_28__N_1411[11]), .S1(multOut_28__N_1411[12])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_4 (.A0(s_mult_29s_25s_0_7_13), .A1(s_mult_29s_25s_0_7_14), 
           .B0(s_mult_29s_25s_0_8_13), .B1(s_mult_29s_25s_0_8_14), .CI(co_mult_29s_25s_0_10_3), 
           .COUT(co_mult_29s_25s_0_10_4), .S0(multOut_28__N_1411[13]), .S1(multOut_28__N_1411[14])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_5 (.A0(s_mult_29s_25s_0_7_15), .A1(s_mult_29s_25s_0_7_16), 
           .B0(s_mult_29s_25s_0_8_15), .B1(s_mult_29s_25s_0_8_16), .CI(co_mult_29s_25s_0_10_4), 
           .COUT(co_mult_29s_25s_0_10_5), .S0(multOut_28__N_1411[15]), .S1(s_mult_29s_25s_0_10_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_6 (.A0(s_mult_29s_25s_0_7_17), .A1(s_mult_29s_25s_0_7_18), 
           .B0(s_mult_29s_25s_0_8_17), .B1(s_mult_29s_25s_0_8_18), .CI(co_mult_29s_25s_0_10_5), 
           .COUT(co_mult_29s_25s_0_10_6), .S0(s_mult_29s_25s_0_10_17), .S1(s_mult_29s_25s_0_10_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_7 (.A0(s_mult_29s_25s_0_7_19), .A1(s_mult_29s_25s_0_7_20), 
           .B0(s_mult_29s_25s_0_8_19), .B1(s_mult_29s_25s_0_8_20), .CI(co_mult_29s_25s_0_10_6), 
           .COUT(co_mult_29s_25s_0_10_7), .S0(s_mult_29s_25s_0_10_19), .S1(s_mult_29s_25s_0_10_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_8 (.A0(s_mult_29s_25s_0_7_21), .A1(s_mult_29s_25s_0_7_22), 
           .B0(s_mult_29s_25s_0_8_21), .B1(s_mult_29s_25s_0_8_22), .CI(co_mult_29s_25s_0_10_7), 
           .COUT(co_mult_29s_25s_0_10_8), .S0(s_mult_29s_25s_0_10_21), .S1(s_mult_29s_25s_0_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_9 (.A0(s_mult_29s_25s_0_7_23), .A1(s_mult_29s_25s_0_7_24), 
           .B0(s_mult_29s_25s_0_8_23), .B1(s_mult_29s_25s_0_8_24), .CI(co_mult_29s_25s_0_10_8), 
           .COUT(co_mult_29s_25s_0_10_9), .S0(s_mult_29s_25s_0_10_23), .S1(s_mult_29s_25s_0_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_10 (.A0(s_mult_29s_25s_0_7_25), .A1(s_mult_29s_25s_0_7_26), 
           .B0(s_mult_29s_25s_0_8_25), .B1(s_mult_29s_25s_0_8_26), .CI(co_mult_29s_25s_0_10_9), 
           .COUT(co_mult_29s_25s_0_10_10), .S0(s_mult_29s_25s_0_10_25), 
           .S1(s_mult_29s_25s_0_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_11 (.A0(s_mult_29s_25s_0_7_27), .A1(s_mult_29s_25s_0_7_28), 
           .B0(s_mult_29s_25s_0_8_27), .B1(s_mult_29s_25s_0_8_28), .CI(co_mult_29s_25s_0_10_10), 
           .S0(s_mult_29s_25s_0_10_27), .S1(s_mult_29s_25s_0_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i10_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[9] ), 
         .D(subIn2_24__N_1534[9]), .Z(subIn2_24__N_1348[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i9_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[8] ), 
         .D(subIn2_24__N_1534[8]), .Z(subIn2_24__N_1348[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i9_3_lut_4_lut.init = 16'hfb40;
    CCU2D sub_16_rep_3_add_2_3 (.A0(n2353[1]), .B0(n4427), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[2]), .B1(n4426), .C1(GND_net), .D1(GND_net), 
          .CIN(n18657), .COUT(n18658), .S0(n4474), .S1(n4473));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_3.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_3.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_3.INJECT1_1 = "NO";
    FADD2B Cadd_mult_29s_25s_0_11_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_9_24), 
           .B0(GND_net), .B1(s_mult_29s_25s_0_6_24), .CI(GND_net), .COUT(co_mult_29s_25s_0_11_1), 
           .S1(s_mult_29s_25s_0_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_2 (.A0(s_mult_29s_25s_0_9_25), .A1(s_mult_29s_25s_0_9_26), 
           .B0(s_mult_29s_25s_0_6_25), .B1(s_mult_29s_25s_0_6_26), .CI(co_mult_29s_25s_0_11_1), 
           .COUT(co_mult_29s_25s_0_11_2), .S0(s_mult_29s_25s_0_11_25), .S1(s_mult_29s_25s_0_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_3 (.A0(s_mult_29s_25s_0_9_27), .A1(s_mult_29s_25s_0_9_28), 
           .B0(s_mult_29s_25s_0_6_27), .B1(s_mult_29s_25s_0_6_28), .CI(co_mult_29s_25s_0_11_2), 
           .S0(s_mult_29s_25s_0_11_27), .S1(s_mult_29s_25s_0_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i8_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[7] ), 
         .D(subIn2_24__N_1534[7]), .Z(subIn2_24__N_1348[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i8_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_t_mult_29s_25s_0_12_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_10_16), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_8_16), .CI(GND_net), .COUT(co_t_mult_29s_25s_0_12_1), 
           .S1(multOut_28__N_1411[16])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_2 (.A0(s_mult_29s_25s_0_10_17), .A1(s_mult_29s_25s_0_10_18), 
           .B0(mult_29s_25s_0_pp_8_17), .B1(s_mult_29s_25s_0_4_18), .CI(co_t_mult_29s_25s_0_12_1), 
           .COUT(co_t_mult_29s_25s_0_12_2), .S0(multOut_28__N_1411[17]), 
           .S1(multOut_28__N_1411[18])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_3 (.A0(s_mult_29s_25s_0_10_19), .A1(s_mult_29s_25s_0_10_20), 
           .B0(s_mult_29s_25s_0_4_19), .B1(s_mult_29s_25s_0_9_20), .CI(co_t_mult_29s_25s_0_12_2), 
           .COUT(co_t_mult_29s_25s_0_12_3), .S0(multOut_28__N_1411[19]), 
           .S1(multOut_28__N_1411[20])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_4 (.A0(s_mult_29s_25s_0_10_21), .A1(s_mult_29s_25s_0_10_22), 
           .B0(s_mult_29s_25s_0_9_21), .B1(s_mult_29s_25s_0_9_22), .CI(co_t_mult_29s_25s_0_12_3), 
           .COUT(co_t_mult_29s_25s_0_12_4), .S0(multOut_28__N_1411[21]), 
           .S1(multOut_28__N_1411[22])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_5 (.A0(s_mult_29s_25s_0_10_23), .A1(s_mult_29s_25s_0_10_24), 
           .B0(s_mult_29s_25s_0_9_23), .B1(s_mult_29s_25s_0_11_24), .CI(co_t_mult_29s_25s_0_12_4), 
           .COUT(co_t_mult_29s_25s_0_12_5), .S0(multOut_28__N_1411[23]), 
           .S1(multOut_28__N_1411[24])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_6 (.A0(s_mult_29s_25s_0_10_25), .A1(s_mult_29s_25s_0_10_26), 
           .B0(s_mult_29s_25s_0_11_25), .B1(s_mult_29s_25s_0_11_26), .CI(co_t_mult_29s_25s_0_12_5), 
           .COUT(co_t_mult_29s_25s_0_12_6), .S0(multOut_28__N_1411[25]), 
           .S1(multOut_28__N_1411[26])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_7 (.A0(s_mult_29s_25s_0_10_27), .A1(s_mult_29s_25s_0_10_28), 
           .B0(s_mult_29s_25s_0_11_27), .B1(s_mult_29s_25s_0_11_28), .CI(co_t_mult_29s_25s_0_12_6), 
           .S0(multOut_28__N_1411[27]), .S1(multOut_28__N_1411[28])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 mux_135_i13_4_lut (.A(backOut2[12]), .B(backOut3[12]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i13_4_lut.init = 16'h0aca;
    MULT2 mult_29s_25s_0_mult_0_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(n21660), .B2(GND_net), .B3(n21660), 
          .CI(mult_29s_25s_0_cin_lr_0), .CO(mco), .P0(multOut_28__N_1411[1]), 
          .P1(mult_29s_25s_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(n21660), .B2(GND_net), .B3(n21660), 
          .CI(mco), .CO(mco_1), .P0(mult_29s_25s_0_pp_0_3), .P1(mult_29s_25s_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(n21660), .B2(GND_net), .B3(n21660), 
          .CI(mco_1), .CO(mco_2), .P0(mult_29s_25s_0_pp_0_5), .P1(mult_29s_25s_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(n21660), .B2(GND_net), .B3(n21660), 
          .CI(mco_2), .CO(mco_3), .P0(mult_29s_25s_0_pp_0_7), .P1(mult_29s_25s_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_3), .CO(mco_4), .P0(mult_29s_25s_0_pp_0_9), 
          .P1(mult_29s_25s_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_4), .CO(mco_5), .P0(mult_29s_25s_0_pp_0_11), 
          .P1(mult_29s_25s_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_5), .CO(mco_6), .P0(mult_29s_25s_0_pp_0_13), 
          .P1(mult_29s_25s_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_6), .CO(mco_7), .P0(mult_29s_25s_0_pp_0_15), 
          .P1(mult_29s_25s_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_7), .CO(mco_8), .P0(mult_29s_25s_0_pp_0_17), 
          .P1(mult_29s_25s_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_8), .CO(mco_9), .P0(mult_29s_25s_0_pp_0_19), 
          .P1(mult_29s_25s_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_9), .CO(mco_10), .P0(mult_29s_25s_0_pp_0_21), 
          .P1(mult_29s_25s_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_10), .CO(mco_11), .P0(mult_29s_25s_0_pp_0_23), 
          .P1(mult_29s_25s_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_11), .CO(mco_12), .P0(mult_29s_25s_0_pp_0_25), 
          .P1(mult_29s_25s_0_pp_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_13 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(n21660), .B2(GND_net), 
          .B3(n21660), .CI(mco_12), .P0(mult_29s_25s_0_pp_0_27), .P1(mult_29s_25s_0_pp_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mult_29s_25s_0_cin_lr_2), .CO(mco_14), 
          .P0(mult_29s_25s_0_pp_1_3), .P1(mult_29s_25s_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_14), .CO(mco_15), .P0(mult_29s_25s_0_pp_1_5), 
          .P1(mult_29s_25s_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_15), .CO(mco_16), .P0(mult_29s_25s_0_pp_1_7), 
          .P1(mult_29s_25s_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_16), .CO(mco_17), .P0(mult_29s_25s_0_pp_1_9), 
          .P1(mult_29s_25s_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_17), .CO(mco_18), .P0(mult_29s_25s_0_pp_1_11), 
          .P1(mult_29s_25s_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_18), .CO(mco_19), .P0(mult_29s_25s_0_pp_1_13), 
          .P1(mult_29s_25s_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_19), .CO(mco_20), .P0(mult_29s_25s_0_pp_1_15), 
          .P1(mult_29s_25s_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_20), .CO(mco_21), .P0(mult_29s_25s_0_pp_1_17), 
          .P1(mult_29s_25s_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_21), .CO(mco_22), .P0(mult_29s_25s_0_pp_1_19), 
          .P1(mult_29s_25s_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_22), .CO(mco_23), .P0(mult_29s_25s_0_pp_1_21), 
          .P1(mult_29s_25s_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_23), .CO(mco_24), .P0(mult_29s_25s_0_pp_1_23), 
          .P1(mult_29s_25s_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_24), .CO(mco_25), .P0(mult_29s_25s_0_pp_1_25), 
          .P1(mult_29s_25s_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[2]), .B2(GND_net), 
          .B3(multIn2[2]), .CI(mco_25), .P0(mult_29s_25s_0_pp_1_27), .P1(mult_29s_25s_0_pp_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mult_29s_25s_0_cin_lr_4), .CO(mco_28), 
          .P0(mult_29s_25s_0_pp_2_5), .P1(mult_29s_25s_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_28), .CO(mco_29), .P0(mult_29s_25s_0_pp_2_7), 
          .P1(mult_29s_25s_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_29), .CO(mco_30), .P0(mult_29s_25s_0_pp_2_9), 
          .P1(mult_29s_25s_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_30), .CO(mco_31), .P0(mult_29s_25s_0_pp_2_11), 
          .P1(mult_29s_25s_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_31), .CO(mco_32), .P0(mult_29s_25s_0_pp_2_13), 
          .P1(mult_29s_25s_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_32), .CO(mco_33), .P0(mult_29s_25s_0_pp_2_15), 
          .P1(mult_29s_25s_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_33), .CO(mco_34), .P0(mult_29s_25s_0_pp_2_17), 
          .P1(mult_29s_25s_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_34), .CO(mco_35), .P0(mult_29s_25s_0_pp_2_19), 
          .P1(mult_29s_25s_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_35), .CO(mco_36), .P0(mult_29s_25s_0_pp_2_21), 
          .P1(mult_29s_25s_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_36), .CO(mco_37), .P0(mult_29s_25s_0_pp_2_23), 
          .P1(mult_29s_25s_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_37), .CO(mco_38), .P0(mult_29s_25s_0_pp_2_25), 
          .P1(mult_29s_25s_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[2]), .B1(multIn2[8]), .B2(multIn2[2]), 
          .B3(multIn2[8]), .CI(mco_38), .P0(mult_29s_25s_0_pp_2_27), .P1(mult_29s_25s_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mult_29s_25s_0_cin_lr_6), .CO(mco_42), 
          .P0(mult_29s_25s_0_pp_3_7), .P1(mult_29s_25s_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_42), .CO(mco_43), .P0(mult_29s_25s_0_pp_3_9), 
          .P1(mult_29s_25s_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_43), .CO(mco_44), .P0(mult_29s_25s_0_pp_3_11), 
          .P1(mult_29s_25s_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_44), .CO(mco_45), .P0(mult_29s_25s_0_pp_3_13), 
          .P1(mult_29s_25s_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_45), .CO(mco_46), .P0(mult_29s_25s_0_pp_3_15), 
          .P1(mult_29s_25s_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_46), .CO(mco_47), .P0(mult_29s_25s_0_pp_3_17), 
          .P1(mult_29s_25s_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_47), .CO(mco_48), .P0(mult_29s_25s_0_pp_3_19), 
          .P1(mult_29s_25s_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_48), .CO(mco_49), .P0(mult_29s_25s_0_pp_3_21), 
          .P1(mult_29s_25s_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_49), .CO(mco_50), .P0(mult_29s_25s_0_pp_3_23), 
          .P1(mult_29s_25s_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_50), .CO(mco_51), .P0(mult_29s_25s_0_pp_3_25), 
          .P1(mult_29s_25s_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[8]), .B1(multIn2[8]), .B2(multIn2[8]), 
          .B3(multIn2[8]), .CI(mco_51), .P0(mult_29s_25s_0_pp_3_27), .P1(mult_29s_25s_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mult_29s_25s_0_cin_lr_8), .CO(mco_56), 
          .P0(mult_29s_25s_0_pp_4_9), .P1(mult_29s_25s_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_56), .CO(mco_57), .P0(mult_29s_25s_0_pp_4_11), 
          .P1(mult_29s_25s_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_57), .CO(mco_58), .P0(mult_29s_25s_0_pp_4_13), 
          .P1(mult_29s_25s_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_58), .CO(mco_59), .P0(mult_29s_25s_0_pp_4_15), 
          .P1(mult_29s_25s_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_59), .CO(mco_60), .P0(mult_29s_25s_0_pp_4_17), 
          .P1(mult_29s_25s_0_pp_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_60), .CO(mco_61), .P0(mult_29s_25s_0_pp_4_19), 
          .P1(mult_29s_25s_0_pp_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_61), .CO(mco_62), .P0(mult_29s_25s_0_pp_4_21), 
          .P1(mult_29s_25s_0_pp_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_62), .CO(mco_63), .P0(mult_29s_25s_0_pp_4_23), 
          .P1(mult_29s_25s_0_pp_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_63), .CO(mco_64), .P0(mult_29s_25s_0_pp_4_25), 
          .P1(mult_29s_25s_0_pp_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[10]), .B1(multIn2[8]), .B2(multIn2[10]), 
          .B3(multIn2[8]), .CI(mco_64), .P0(mult_29s_25s_0_pp_4_27), .P1(mult_29s_25s_0_pp_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i4_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[3] ), 
         .D(subIn2_24__N_1534[3]), .Z(subIn2_24__N_1348[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i4_3_lut_4_lut.init = 16'hfb40;
    MULT2 mult_29s_25s_0_mult_10_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mult_29s_25s_0_cin_lr_10), .CO(mco_70), 
          .P0(mult_29s_25s_0_pp_5_11), .P1(mult_29s_25s_0_pp_5_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_70), .CO(mco_71), .P0(mult_29s_25s_0_pp_5_13), 
          .P1(mult_29s_25s_0_pp_5_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_71), .CO(mco_72), .P0(mult_29s_25s_0_pp_5_15), 
          .P1(mult_29s_25s_0_pp_5_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_72), .CO(mco_73), .P0(mult_29s_25s_0_pp_5_17), 
          .P1(mult_29s_25s_0_pp_5_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_73), .CO(mco_74), .P0(mult_29s_25s_0_pp_5_19), 
          .P1(mult_29s_25s_0_pp_5_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_74), .CO(mco_75), .P0(mult_29s_25s_0_pp_5_21), 
          .P1(mult_29s_25s_0_pp_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_75), .CO(mco_76), .P0(mult_29s_25s_0_pp_5_23), 
          .P1(mult_29s_25s_0_pp_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_76), .CO(mco_77), .P0(mult_29s_25s_0_pp_5_25), 
          .P1(mult_29s_25s_0_pp_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(multIn2[10]), .B2(GND_net), 
          .B3(multIn2[10]), .CI(mco_77), .P0(mult_29s_25s_0_pp_5_27), 
          .P1(mult_29s_25s_0_pp_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i20_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[19] ), 
         .D(\speed_avg_m2[19] ), .Z(subIn2_24__N_1348[19])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3326_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m2[9]), .Z(n5821)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3326_3_lut_4_lut.init = 16'hfd20;
    MULT2 mult_29s_25s_0_mult_12_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_12), .CO(mco_84), .P0(mult_29s_25s_0_pp_6_13), 
          .P1(mult_29s_25s_0_pp_6_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_84), .CO(mco_85), .P0(mult_29s_25s_0_pp_6_15), 
          .P1(mult_29s_25s_0_pp_6_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_85), .CO(mco_86), .P0(mult_29s_25s_0_pp_6_17), 
          .P1(mult_29s_25s_0_pp_6_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_86), .CO(mco_87), .P0(mult_29s_25s_0_pp_6_19), 
          .P1(mult_29s_25s_0_pp_6_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_87), .CO(mco_88), .P0(mult_29s_25s_0_pp_6_21), 
          .P1(mult_29s_25s_0_pp_6_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_88), .CO(mco_89), .P0(mult_29s_25s_0_pp_6_23), 
          .P1(mult_29s_25s_0_pp_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_89), .CO(mco_90), .P0(mult_29s_25s_0_pp_6_25), 
          .P1(mult_29s_25s_0_pp_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_90), .P0(mult_29s_25s_0_pp_6_27), .P1(mult_29s_25s_0_pp_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_14), .CO(mco_98), .P0(mult_29s_25s_0_pp_7_15), 
          .P1(mult_29s_25s_0_pp_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_98), .CO(mco_99), .P0(mult_29s_25s_0_pp_7_17), 
          .P1(mult_29s_25s_0_pp_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_99), .CO(mco_100), .P0(mult_29s_25s_0_pp_7_19), 
          .P1(mult_29s_25s_0_pp_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_100), .CO(mco_101), .P0(mult_29s_25s_0_pp_7_21), 
          .P1(mult_29s_25s_0_pp_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_101), .CO(mco_102), .P0(mult_29s_25s_0_pp_7_23), 
          .P1(mult_29s_25s_0_pp_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_102), .CO(mco_103), .P0(mult_29s_25s_0_pp_7_25), 
          .P1(mult_29s_25s_0_pp_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_103), .P0(mult_29s_25s_0_pp_7_27), .P1(mult_29s_25s_0_pp_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_16), .CO(mco_112), .P0(mult_29s_25s_0_pp_8_17), 
          .P1(mult_29s_25s_0_pp_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_112), .CO(mco_113), .P0(mult_29s_25s_0_pp_8_19), 
          .P1(mult_29s_25s_0_pp_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_113), .CO(mco_114), .P0(mult_29s_25s_0_pp_8_21), 
          .P1(mult_29s_25s_0_pp_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_114), .CO(mco_115), .P0(mult_29s_25s_0_pp_8_23), 
          .P1(mult_29s_25s_0_pp_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_115), .CO(mco_116), .P0(mult_29s_25s_0_pp_8_25), 
          .P1(mult_29s_25s_0_pp_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_116), .P0(mult_29s_25s_0_pp_8_27), .P1(mult_29s_25s_0_pp_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i19_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[18] ), 
         .D(\speed_avg_m2[18] ), .Z(subIn2_24__N_1348[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i18_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[17] ), 
         .D(\speed_avg_m2[17] ), .Z(subIn2_24__N_1348[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i18_3_lut_4_lut.init = 16'hfb40;
    MULT2 mult_29s_25s_0_mult_18_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_18), .CO(mco_126), .P0(mult_29s_25s_0_pp_9_19), 
          .P1(mult_29s_25s_0_pp_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_126), .CO(mco_127), .P0(mult_29s_25s_0_pp_9_21), 
          .P1(mult_29s_25s_0_pp_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_127), .CO(mco_128), .P0(mult_29s_25s_0_pp_9_23), 
          .P1(mult_29s_25s_0_pp_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_128), .CO(mco_129), .P0(mult_29s_25s_0_pp_9_25), 
          .P1(mult_29s_25s_0_pp_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_129), .P0(mult_29s_25s_0_pp_9_27), .P1(mult_29s_25s_0_pp_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_20), .CO(mco_140), .P0(mult_29s_25s_0_pp_10_21), 
          .P1(mult_29s_25s_0_pp_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_140), .CO(mco_141), .P0(mult_29s_25s_0_pp_10_23), 
          .P1(mult_29s_25s_0_pp_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_141), .CO(mco_142), .P0(mult_29s_25s_0_pp_10_25), 
          .P1(mult_29s_25s_0_pp_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_142), .P0(mult_29s_25s_0_pp_10_27), .P1(mult_29s_25s_0_pp_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i17_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[16] ), 
         .D(\speed_avg_m2[16] ), .Z(subIn2_24__N_1348[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i17_3_lut_4_lut.init = 16'hfb40;
    PFUMX i17825 (.BLUT(n22420), .ALUT(n22421), .C0(ss[1]), .Z(n16309));
    LUT4 subIn2_24__I_25_i16_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[15] ), 
         .D(\speed_avg_m2[15] ), .Z(subIn2_24__N_1348[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i16_3_lut_4_lut.init = 16'hfb40;
    MULT2 mult_29s_25s_0_mult_22_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_22), .CO(mco_154), .P0(mult_29s_25s_0_pp_11_23), 
          .P1(mult_29s_25s_0_pp_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_154), .CO(mco_155), .P0(mult_29s_25s_0_pp_11_25), 
          .P1(mult_29s_25s_0_pp_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_155), .P0(mult_29s_25s_0_pp_11_27), .P1(mult_29s_25s_0_pp_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 mux_135_i14_4_lut (.A(backOut2[13]), .B(backOut3[13]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i14_4_lut.init = 16'h0aca;
    LUT4 subIn2_24__I_25_i15_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[14] ), 
         .D(\speed_avg_m2[14] ), .Z(subIn2_24__N_1348[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17498_2_lut_rep_317_2_lut_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), 
         .C(n42), .D(n16309), .Z(n21630)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (C+(D)))) */ ;
    defparam i17498_2_lut_rep_317_2_lut_3_lut_4_lut.init = 16'h222f;
    LUT4 subIn2_24__I_25_i14_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[13] ), 
         .D(\speed_avg_m2[13] ), .Z(subIn2_24__N_1348[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i12_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[11] ), 
         .D(\speed_avg_m2[11] ), .Z(subIn2_24__N_1348[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i12_3_lut_4_lut.init = 16'hfb40;
    FADD2B mult_29s_25s_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i13240_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[3]), 
         .D(ss[1]), .Z(intgOut3_28__N_1058[3])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13240_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 subIn2_24__I_25_i11_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[10] ), 
         .D(\speed_avg_m2[10] ), .Z(subIn2_24__N_1348[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_189_i10_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[9]), 
         .Z(intgOut0_28__N_1627[9])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i10_3_lut_3_lut.init = 16'hbaba;
    LUT4 i13239_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[4]), 
         .D(ss[1]), .Z(intgOut3_28__N_1058[4])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13239_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 subIn2_24__I_25_i7_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[6] ), 
         .D(\speed_avg_m2[6] ), .Z(subIn2_24__N_1348[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i6_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[5] ), 
         .D(\speed_avg_m2[5] ), .Z(subIn2_24__N_1348[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i5_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[4] ), 
         .D(\speed_avg_m2[4] ), .Z(subIn2_24__N_1348[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13136_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[0]), 
         .D(ss[1]), .Z(intgOut2_28__N_1029[0])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13136_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_135_i15_4_lut (.A(backOut2[14]), .B(backOut3[14]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i15_4_lut.init = 16'h0aca;
    LUT4 i3023_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m2[0]), .Z(n5518)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3023_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_64 (.A(n21725), .B(n19907), .C(n22440), .D(n21697), 
         .Z(clk_N_875_enable_220)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_64.init = 16'hc0c8;
    LUT4 subIn2_24__I_25_i3_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[2] ), 
         .D(\speed_avg_m2[2] ), .Z(subIn2_24__N_1348[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_adj_65 (.A(n21725), .B(n19907), .C(n22440), .D(n21726), 
         .Z(clk_N_875_enable_248)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_65.init = 16'hc8c0;
    LUT4 subIn2_24__I_25_i2_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[1] ), 
         .D(\speed_avg_m2[1] ), .Z(subIn2_24__N_1348[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i1_3_lut_4_lut (.A(ss[2]), .B(n21688), .C(\speed_avg_m1[0] ), 
         .D(\speed_avg_m2[0] ), .Z(subIn2_24__N_1348[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i17541_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut_4_lut (.A(n21729), .B(ss[0]), 
         .C(ss[2]), .D(ss[1]), .Z(n20645)) /* synthesis lut_function=(!(A+(B (C (D))+!B !(C+(D))))) */ ;
    defparam i17541_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut_4_lut.init = 16'h1554;
    LUT4 i17475_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21686), .D(n22424), .Z(n20372)) /* synthesis lut_function=(!((B (C (D))+!B (D))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam i17475_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h08aa;
    LUT4 i3310_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m2[1]), .Z(n5805)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3310_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i16_4_lut (.A(backOut2[15]), .B(backOut3[15]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i16_4_lut.init = 16'h0aca;
    LUT4 i3312_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m2[2]), .Z(n5807)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3312_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3314_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m2[3]), .Z(n5809)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3314_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3316_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m2[4]), .Z(n5811)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3316_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i17_4_lut (.A(backOut2[16]), .B(backOut3[16]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i17_4_lut.init = 16'h0aca;
    LUT4 i3318_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m2[5]), .Z(n5813)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3318_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3320_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m2[6]), .Z(n5815)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3320_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3322_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m2[7]), .Z(n5817)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3322_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3324_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m2[8]), .Z(n5819)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3324_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX backOut0_i0_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_72), 
            .CK(clk_N_875), .Q(backOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i1.GSR = "DISABLED";
    FD1S3AX multOut_i1 (.D(multOut_28__N_1411[1]), .CK(clk_N_875), .Q(multOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i1.GSR = "ENABLED";
    LUT4 mux_189_i21_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[20]), 
         .Z(intgOut0_28__N_1627[20])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i21_3_lut_3_lut.init = 16'hbaba;
    CCU2D sub_16_rep_3_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[0]), .B1(n4428), .C1(GND_net), .D1(GND_net), 
          .COUT(n18657), .S1(n4475));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_1.INIT0 = 16'h0000;
    defparam sub_16_rep_3_add_2_1.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_1.INJECT1_1 = "NO";
    CCU2D add_15377_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18656), 
          .S0(n3636));
    defparam add_15377_cout.INIT0 = 16'h0000;
    defparam add_15377_cout.INIT1 = 16'h0000;
    defparam add_15377_cout.INJECT1_0 = "NO";
    defparam add_15377_cout.INJECT1_1 = "NO";
    LUT4 i3328_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m2[10]), .Z(n5823)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3328_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15377_20 (.A0(speed_set_m1[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18655), .COUT(n18656));
    defparam add_15377_20.INIT0 = 16'h5aaa;
    defparam add_15377_20.INIT1 = 16'h0aaa;
    defparam add_15377_20.INJECT1_0 = "NO";
    defparam add_15377_20.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(ss[3]), .B(n22425), .C(ss[0]), .D(ss[1]), .Z(subIn1_24__N_1342)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C (D)+!C !(D))))) */ ;
    defparam i2_4_lut.init = 16'h0130;
    CCU2D add_15377_18 (.A0(speed_set_m1[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18654), .COUT(n18655));
    defparam add_15377_18.INIT0 = 16'h5aaa;
    defparam add_15377_18.INIT1 = 16'h5aaa;
    defparam add_15377_18.INJECT1_0 = "NO";
    defparam add_15377_18.INJECT1_1 = "NO";
    CCU2D add_15377_16 (.A0(speed_set_m1[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18653), .COUT(n18654));
    defparam add_15377_16.INIT0 = 16'h5aaa;
    defparam add_15377_16.INIT1 = 16'h5aaa;
    defparam add_15377_16.INJECT1_0 = "NO";
    defparam add_15377_16.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_66 (.A(n21635), .B(n22418), .C(n21634), .D(n56), 
         .Z(n16073)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i2_4_lut_adj_66.init = 16'hfbfa;
    CCU2D add_15377_14 (.A0(speed_set_m1[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18652), .COUT(n18653));
    defparam add_15377_14.INIT0 = 16'h5555;
    defparam add_15377_14.INIT1 = 16'h5aaa;
    defparam add_15377_14.INJECT1_0 = "NO";
    defparam add_15377_14.INJECT1_1 = "NO";
    CCU2D add_15377_12 (.A0(speed_set_m1[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18651), .COUT(n18652));
    defparam add_15377_12.INIT0 = 16'h5aaa;
    defparam add_15377_12.INIT1 = 16'h5aaa;
    defparam add_15377_12.INJECT1_0 = "NO";
    defparam add_15377_12.INJECT1_1 = "NO";
    LUT4 i3330_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m2[11]), .Z(n5825)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3330_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15370_29 (.A0(addOut[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18768), 
          .S1(n3844));
    defparam add_15370_29.INIT0 = 16'h5aaa;
    defparam add_15370_29.INIT1 = 16'h0000;
    defparam add_15370_29.INJECT1_0 = "NO";
    defparam add_15370_29.INJECT1_1 = "NO";
    CCU2D add_15370_27 (.A0(addOut[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18767), .COUT(n18768));
    defparam add_15370_27.INIT0 = 16'h0aaa;
    defparam add_15370_27.INIT1 = 16'h0aaa;
    defparam add_15370_27.INJECT1_0 = "NO";
    defparam add_15370_27.INJECT1_1 = "NO";
    CCU2D add_15370_25 (.A0(addOut[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18766), .COUT(n18767));
    defparam add_15370_25.INIT0 = 16'h0aaa;
    defparam add_15370_25.INIT1 = 16'h0aaa;
    defparam add_15370_25.INJECT1_0 = "NO";
    defparam add_15370_25.INJECT1_1 = "NO";
    LUT4 i13134_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[1]), 
         .D(ss[1]), .Z(intgOut2_28__N_1029[1])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13134_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i13133_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[2]), 
         .D(ss[1]), .Z(intgOut2_28__N_1029[2])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13133_2_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D add_15377_10 (.A0(speed_set_m1[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18650), .COUT(n18651));
    defparam add_15377_10.INIT0 = 16'h5555;
    defparam add_15377_10.INIT1 = 16'h5555;
    defparam add_15377_10.INJECT1_0 = "NO";
    defparam add_15377_10.INJECT1_1 = "NO";
    LUT4 i13130_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[3]), 
         .D(ss[1]), .Z(intgOut2_28__N_1029[3])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13130_2_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D add_15370_23 (.A0(addOut[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18765), .COUT(n18766));
    defparam add_15370_23.INIT0 = 16'h0aaa;
    defparam add_15370_23.INIT1 = 16'h0aaa;
    defparam add_15370_23.INJECT1_0 = "NO";
    defparam add_15370_23.INJECT1_1 = "NO";
    LUT4 i13129_2_lut_3_lut_4_lut (.A(n21687), .B(n21628), .C(addOut[4]), 
         .D(ss[1]), .Z(intgOut2_28__N_1029[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13129_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i3332_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m2[12]), .Z(n5827)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3332_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2_4_lut_adj_67 (.A(n21666), .B(n22424), .C(n21723), .D(n6), 
         .Z(n15564)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i2_4_lut_adj_67.init = 16'ha888;
    LUT4 i3334_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m2[13]), .Z(n5829)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3334_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i18_4_lut (.A(backOut2[17]), .B(backOut3[17]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i18_4_lut.init = 16'h0aca;
    CCU2D add_15377_8 (.A0(speed_set_m1[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18649), .COUT(n18650));
    defparam add_15377_8.INIT0 = 16'h5aaa;
    defparam add_15377_8.INIT1 = 16'h5555;
    defparam add_15377_8.INJECT1_0 = "NO";
    defparam add_15377_8.INJECT1_1 = "NO";
    LUT4 i3336_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m2[14]), .Z(n5831)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3336_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15370_21 (.A0(addOut[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18764), .COUT(n18765));
    defparam add_15370_21.INIT0 = 16'hf555;
    defparam add_15370_21.INIT1 = 16'h0aaa;
    defparam add_15370_21.INJECT1_0 = "NO";
    defparam add_15370_21.INJECT1_1 = "NO";
    LUT4 i3338_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m2[15]), .Z(n5833)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3338_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15370_19 (.A0(addOut[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18763), .COUT(n18764));
    defparam add_15370_19.INIT0 = 16'hf555;
    defparam add_15370_19.INIT1 = 16'h0aaa;
    defparam add_15370_19.INJECT1_0 = "NO";
    defparam add_15370_19.INJECT1_1 = "NO";
    CCU2D add_15370_17 (.A0(addOut[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18762), .COUT(n18763));
    defparam add_15370_17.INIT0 = 16'h0aaa;
    defparam add_15370_17.INIT1 = 16'hf555;
    defparam add_15370_17.INJECT1_0 = "NO";
    defparam add_15370_17.INJECT1_1 = "NO";
    CCU2D add_15377_6 (.A0(speed_set_m1[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18648), .COUT(n18649));
    defparam add_15377_6.INIT0 = 16'h5aaa;
    defparam add_15377_6.INIT1 = 16'h5aaa;
    defparam add_15377_6.INJECT1_0 = "NO";
    defparam add_15377_6.INJECT1_1 = "NO";
    CCU2D add_15377_4 (.A0(speed_set_m1[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18647), .COUT(n18648));
    defparam add_15377_4.INIT0 = 16'h5555;
    defparam add_15377_4.INIT1 = 16'h5aaa;
    defparam add_15377_4.INJECT1_0 = "NO";
    defparam add_15377_4.INJECT1_1 = "NO";
    CCU2D add_15370_15 (.A0(addOut[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18761), .COUT(n18762));
    defparam add_15370_15.INIT0 = 16'hf555;
    defparam add_15370_15.INIT1 = 16'hf555;
    defparam add_15370_15.INJECT1_0 = "NO";
    defparam add_15370_15.INJECT1_1 = "NO";
    CCU2D add_15377_2 (.A0(speed_set_m1[1]), .B0(speed_set_m1[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18647));
    defparam add_15377_2.INIT0 = 16'h1000;
    defparam add_15377_2.INIT1 = 16'h5555;
    defparam add_15377_2.INJECT1_0 = "NO";
    defparam add_15377_2.INJECT1_1 = "NO";
    CCU2D add_15370_13 (.A0(addOut[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18760), .COUT(n18761));
    defparam add_15370_13.INIT0 = 16'h0aaa;
    defparam add_15370_13.INIT1 = 16'hf555;
    defparam add_15370_13.INJECT1_0 = "NO";
    defparam add_15370_13.INJECT1_1 = "NO";
    CCU2D add_15370_11 (.A0(addOut[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18759), .COUT(n18760));
    defparam add_15370_11.INIT0 = 16'h0aaa;
    defparam add_15370_11.INIT1 = 16'h0aaa;
    defparam add_15370_11.INJECT1_0 = "NO";
    defparam add_15370_11.INJECT1_1 = "NO";
    CCU2D add_15378_17 (.A0(speed_set_m1[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18646), .S1(n3612));
    defparam add_15378_17.INIT0 = 16'h5555;
    defparam add_15378_17.INIT1 = 16'h0000;
    defparam add_15378_17.INJECT1_0 = "NO";
    defparam add_15378_17.INJECT1_1 = "NO";
    CCU2D add_15378_15 (.A0(speed_set_m1[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18645), .COUT(n18646));
    defparam add_15378_15.INIT0 = 16'hf555;
    defparam add_15378_15.INIT1 = 16'hf555;
    defparam add_15378_15.INJECT1_0 = "NO";
    defparam add_15378_15.INJECT1_1 = "NO";
    CCU2D add_15378_13 (.A0(speed_set_m1[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18644), .COUT(n18645));
    defparam add_15378_13.INIT0 = 16'hf555;
    defparam add_15378_13.INIT1 = 16'hf555;
    defparam add_15378_13.INJECT1_0 = "NO";
    defparam add_15378_13.INJECT1_1 = "NO";
    CCU2D add_15370_9 (.A0(addOut[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18758), .COUT(n18759));
    defparam add_15370_9.INIT0 = 16'hf555;
    defparam add_15370_9.INIT1 = 16'hf555;
    defparam add_15370_9.INJECT1_0 = "NO";
    defparam add_15370_9.INJECT1_1 = "NO";
    LUT4 i3340_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m2[16]), .Z(n5835)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3340_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i19_4_lut (.A(backOut2[18]), .B(backOut3[18]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i19_4_lut.init = 16'h0aca;
    LUT4 i3342_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m2[17]), .Z(n5837)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3342_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3344_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m2[18]), .Z(n5839)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3344_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i20_4_lut (.A(backOut2[19]), .B(backOut3[19]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i20_4_lut.init = 16'h0aca;
    LUT4 i3346_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m2[19]), .Z(n5841)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3346_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3350_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m2[20]), .Z(n5845)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3350_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i21_4_lut (.A(backOut2[20]), .B(backOut3[20]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i21_4_lut.init = 16'h0aca;
    CCU2D add_15378_11 (.A0(speed_set_m1[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18643), .COUT(n18644));
    defparam add_15378_11.INIT0 = 16'hf555;
    defparam add_15378_11.INIT1 = 16'hf555;
    defparam add_15378_11.INJECT1_0 = "NO";
    defparam add_15378_11.INJECT1_1 = "NO";
    CCU2D add_15370_7 (.A0(addOut[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18757), .COUT(n18758));
    defparam add_15370_7.INIT0 = 16'hf555;
    defparam add_15370_7.INIT1 = 16'h0aaa;
    defparam add_15370_7.INJECT1_0 = "NO";
    defparam add_15370_7.INJECT1_1 = "NO";
    FD1S3AX multOut_i2 (.D(multOut_28__N_1411[2]), .CK(clk_N_875), .Q(multOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i2.GSR = "ENABLED";
    FD1S3AX multOut_i3 (.D(multOut_28__N_1411[3]), .CK(clk_N_875), .Q(multOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i3.GSR = "ENABLED";
    FD1S3AX multOut_i4 (.D(multOut_28__N_1411[4]), .CK(clk_N_875), .Q(multOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i4.GSR = "ENABLED";
    FD1S3AX multOut_i5 (.D(multOut_28__N_1411[5]), .CK(clk_N_875), .Q(multOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i5.GSR = "ENABLED";
    FD1S3AX multOut_i6 (.D(multOut_28__N_1411[6]), .CK(clk_N_875), .Q(multOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i6.GSR = "ENABLED";
    FD1S3AX multOut_i7 (.D(multOut_28__N_1411[7]), .CK(clk_N_875), .Q(multOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i7.GSR = "ENABLED";
    FD1S3AX multOut_i8 (.D(multOut_28__N_1411[8]), .CK(clk_N_875), .Q(multOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i8.GSR = "ENABLED";
    FD1S3AX multOut_i9 (.D(multOut_28__N_1411[9]), .CK(clk_N_875), .Q(multOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i9.GSR = "ENABLED";
    FD1S3AX multOut_i10 (.D(multOut_28__N_1411[10]), .CK(clk_N_875), .Q(multOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i10.GSR = "ENABLED";
    FD1S3AX multOut_i11 (.D(multOut_28__N_1411[11]), .CK(clk_N_875), .Q(multOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i11.GSR = "ENABLED";
    FD1S3AX multOut_i12 (.D(multOut_28__N_1411[12]), .CK(clk_N_875), .Q(multOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i12.GSR = "ENABLED";
    FD1S3AX multOut_i13 (.D(multOut_28__N_1411[13]), .CK(clk_N_875), .Q(multOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i13.GSR = "ENABLED";
    FD1S3AX multOut_i14 (.D(multOut_28__N_1411[14]), .CK(clk_N_875), .Q(multOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i14.GSR = "ENABLED";
    FD1S3AX multOut_i15 (.D(multOut_28__N_1411[15]), .CK(clk_N_875), .Q(multOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i15.GSR = "ENABLED";
    FD1S3AX multOut_i16 (.D(multOut_28__N_1411[16]), .CK(clk_N_875), .Q(multOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i16.GSR = "ENABLED";
    FD1S3AX multOut_i17 (.D(multOut_28__N_1411[17]), .CK(clk_N_875), .Q(multOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i17.GSR = "ENABLED";
    FD1S3AX multOut_i18 (.D(multOut_28__N_1411[18]), .CK(clk_N_875), .Q(multOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i18.GSR = "ENABLED";
    FD1S3AX multOut_i19 (.D(multOut_28__N_1411[19]), .CK(clk_N_875), .Q(multOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i19.GSR = "ENABLED";
    FD1S3AX multOut_i20 (.D(multOut_28__N_1411[20]), .CK(clk_N_875), .Q(multOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i20.GSR = "ENABLED";
    FD1S3AX multOut_i21 (.D(multOut_28__N_1411[21]), .CK(clk_N_875), .Q(multOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i21.GSR = "ENABLED";
    FD1S3AX multOut_i22 (.D(multOut_28__N_1411[22]), .CK(clk_N_875), .Q(multOut[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i22.GSR = "ENABLED";
    FD1S3AX multOut_i23 (.D(multOut_28__N_1411[23]), .CK(clk_N_875), .Q(multOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i23.GSR = "ENABLED";
    FD1S3AX multOut_i24 (.D(multOut_28__N_1411[24]), .CK(clk_N_875), .Q(multOut[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i24.GSR = "ENABLED";
    FD1S3AX multOut_i25 (.D(multOut_28__N_1411[25]), .CK(clk_N_875), .Q(multOut[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i25.GSR = "ENABLED";
    FD1S3AX multOut_i26 (.D(multOut_28__N_1411[26]), .CK(clk_N_875), .Q(multOut[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i26.GSR = "ENABLED";
    FD1S3AX multOut_i27 (.D(multOut_28__N_1411[27]), .CK(clk_N_875), .Q(multOut[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i27.GSR = "ENABLED";
    FD1S3AX multOut_i28 (.D(multOut_28__N_1411[28]), .CK(clk_N_875), .Q(multOut[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i28.GSR = "ENABLED";
    LUT4 mux_135_i22_4_lut (.A(backOut2[21]), .B(backOut3[21]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i22_4_lut.init = 16'h0aca;
    LUT4 mux_189_i14_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[13]), 
         .Z(intgOut0_28__N_1627[13])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i14_3_lut_3_lut.init = 16'hbaba;
    LUT4 mux_189_i16_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[15]), 
         .Z(intgOut0_28__N_1627[15])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i16_3_lut_3_lut.init = 16'hbaba;
    FD1P3AX intgOut2_i1 (.D(intgOut2_28__N_1029[1]), .SP(clk_N_875_enable_333), 
            .CK(clk_N_875), .Q(intgOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i1.GSR = "ENABLED";
    FD1P3AX intgOut2_i2 (.D(intgOut2_28__N_1029[2]), .SP(clk_N_875_enable_333), 
            .CK(clk_N_875), .Q(intgOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i2.GSR = "ENABLED";
    FD1P3AX intgOut2_i3 (.D(intgOut2_28__N_1029[3]), .SP(clk_N_875_enable_333), 
            .CK(clk_N_875), .Q(intgOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i3.GSR = "ENABLED";
    FD1P3AX intgOut2_i4 (.D(intgOut2_28__N_1029[4]), .SP(clk_N_875_enable_333), 
            .CK(clk_N_875), .Q(intgOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i4.GSR = "ENABLED";
    FD1P3AX intgOut3_i1 (.D(intgOut3_28__N_1058[1]), .SP(clk_N_875_enable_309), 
            .CK(clk_N_875), .Q(intgOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i1.GSR = "ENABLED";
    FD1P3AX intgOut3_i2 (.D(intgOut3_28__N_1058[2]), .SP(clk_N_875_enable_309), 
            .CK(clk_N_875), .Q(intgOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i2.GSR = "ENABLED";
    FD1P3AX intgOut3_i3 (.D(intgOut3_28__N_1058[3]), .SP(clk_N_875_enable_309), 
            .CK(clk_N_875), .Q(intgOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i3.GSR = "ENABLED";
    FD1P3AX intgOut3_i4 (.D(intgOut3_28__N_1058[4]), .SP(clk_N_875_enable_309), 
            .CK(clk_N_875), .Q(intgOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i4.GSR = "ENABLED";
    LUT4 mux_135_i23_4_lut (.A(backOut2[22]), .B(backOut3[22]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i23_4_lut.init = 16'h0aca;
    LUT4 mux_189_i15_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[14]), 
         .Z(intgOut0_28__N_1627[14])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i15_3_lut_3_lut.init = 16'hbaba;
    FD1P3AX Out0_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i1.GSR = "ENABLED";
    FD1P3AX Out0_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i2.GSR = "ENABLED";
    FD1P3AX Out0_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i3.GSR = "ENABLED";
    FD1P3AX Out0_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i4.GSR = "ENABLED";
    FD1P3AX Out0_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i5.GSR = "ENABLED";
    FD1P3AX Out0_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i6.GSR = "ENABLED";
    FD1P3AX Out0_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i7.GSR = "ENABLED";
    FD1P3AX Out0_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i8.GSR = "ENABLED";
    FD1P3AX Out0_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i9.GSR = "ENABLED";
    FD1P3AX Out0_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i10.GSR = "ENABLED";
    FD1P3AX Out0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i11.GSR = "ENABLED";
    FD1P3AX Out0_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i12.GSR = "ENABLED";
    FD1P3AX Out0_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i13.GSR = "ENABLED";
    FD1P3AX Out0_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i14.GSR = "ENABLED";
    FD1P3AX Out0_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i15.GSR = "ENABLED";
    FD1P3AX Out0_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i16.GSR = "ENABLED";
    FD1P3AX Out0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i17.GSR = "ENABLED";
    FD1P3AX Out0_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i18.GSR = "ENABLED";
    FD1P3AX Out0_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i19.GSR = "ENABLED";
    FD1P3AX Out0_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i20.GSR = "ENABLED";
    FD1P3AX Out0_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i21.GSR = "ENABLED";
    FD1P3AX Out0_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i22.GSR = "ENABLED";
    FD1P3AX Out0_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i23.GSR = "ENABLED";
    FD1P3AX Out0_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i24.GSR = "ENABLED";
    FD1P3AX Out0_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i25.GSR = "ENABLED";
    FD1P3AX Out0_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i26.GSR = "ENABLED";
    FD1P3AX Out0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i27.GSR = "ENABLED";
    FD1P3AX Out0_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_108), 
            .CK(clk_N_875), .Q(Out0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i28.GSR = "ENABLED";
    FD1P3AX Out1_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i1.GSR = "ENABLED";
    FD1P3AX Out1_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i2.GSR = "ENABLED";
    FD1P3AX Out1_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i3.GSR = "ENABLED";
    FD1P3AX Out1_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i4.GSR = "ENABLED";
    FD1P3AX Out1_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i5.GSR = "ENABLED";
    FD1P3AX Out1_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i6.GSR = "ENABLED";
    FD1P3AX Out1_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i7.GSR = "ENABLED";
    FD1P3AX Out1_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i8.GSR = "ENABLED";
    FD1P3AX Out1_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i9.GSR = "ENABLED";
    FD1P3AX Out1_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i10.GSR = "ENABLED";
    FD1P3AX Out1_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i11.GSR = "ENABLED";
    FD1P3AX Out1_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i12.GSR = "ENABLED";
    FD1P3AX Out1_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i13.GSR = "ENABLED";
    FD1P3AX Out1_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i14.GSR = "ENABLED";
    FD1P3AX Out1_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i15.GSR = "ENABLED";
    FD1P3AX Out1_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i16.GSR = "ENABLED";
    FD1P3AX Out1_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i17.GSR = "ENABLED";
    FD1P3AX Out1_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i18.GSR = "ENABLED";
    FD1P3AX Out1_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i19.GSR = "ENABLED";
    FD1P3AX Out1_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i20.GSR = "ENABLED";
    FD1P3AX Out1_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i21.GSR = "ENABLED";
    FD1P3AX Out1_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i22.GSR = "ENABLED";
    FD1P3AX Out1_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i23.GSR = "ENABLED";
    FD1P3AX Out1_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i24.GSR = "ENABLED";
    FD1P3AX Out1_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i25.GSR = "ENABLED";
    FD1P3AX Out1_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i26.GSR = "ENABLED";
    FD1P3AX Out1_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i27.GSR = "ENABLED";
    FD1P3AX Out1_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_136), 
            .CK(clk_N_875), .Q(Out1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i28.GSR = "ENABLED";
    FD1P3AX Out2_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i1.GSR = "ENABLED";
    FD1P3AX Out2_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i2.GSR = "ENABLED";
    FD1P3AX Out2_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i3.GSR = "ENABLED";
    FD1P3AX Out2_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i4.GSR = "ENABLED";
    FD1P3AX Out2_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i5.GSR = "ENABLED";
    FD1P3AX Out2_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i6.GSR = "ENABLED";
    FD1P3AX Out2_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i7.GSR = "ENABLED";
    FD1P3AX Out2_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i8.GSR = "ENABLED";
    FD1P3AX Out2_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i9.GSR = "ENABLED";
    FD1P3AX Out2_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i10.GSR = "ENABLED";
    FD1P3AX Out2_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i11.GSR = "ENABLED";
    FD1P3AX Out2_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i12.GSR = "ENABLED";
    FD1P3AX Out2_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i13.GSR = "ENABLED";
    FD1P3AX Out2_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i14.GSR = "ENABLED";
    FD1P3AX Out2_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i15.GSR = "ENABLED";
    FD1P3AX Out2_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i16.GSR = "ENABLED";
    FD1P3AX Out2_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i17.GSR = "ENABLED";
    FD1P3AX Out2_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i18.GSR = "ENABLED";
    FD1P3AX Out2_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i19.GSR = "ENABLED";
    FD1P3AX Out2_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i20.GSR = "ENABLED";
    FD1P3AX Out2_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i21.GSR = "ENABLED";
    FD1P3AX Out2_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i22.GSR = "ENABLED";
    FD1P3AX Out2_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i23.GSR = "ENABLED";
    FD1P3AX Out2_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i24.GSR = "ENABLED";
    FD1P3AX Out2_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i25.GSR = "ENABLED";
    FD1P3AX Out2_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i26.GSR = "ENABLED";
    FD1P3AX Out2_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i27.GSR = "ENABLED";
    FD1P3AX Out2_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_164), 
            .CK(clk_N_875), .Q(Out2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i28.GSR = "ENABLED";
    FD1P3AX Out3_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i1.GSR = "ENABLED";
    FD1P3AX Out3_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i2.GSR = "ENABLED";
    FD1P3AX Out3_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i3.GSR = "ENABLED";
    FD1P3AX Out3_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i4.GSR = "ENABLED";
    FD1P3AX Out3_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i5.GSR = "ENABLED";
    FD1P3AX Out3_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i6.GSR = "ENABLED";
    FD1P3AX Out3_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i7.GSR = "ENABLED";
    FD1P3AX Out3_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i8.GSR = "ENABLED";
    FD1P3AX Out3_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i9.GSR = "ENABLED";
    FD1P3AX Out3_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i10.GSR = "ENABLED";
    FD1P3AX Out3_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i11.GSR = "ENABLED";
    FD1P3AX Out3_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i12.GSR = "ENABLED";
    FD1P3AX Out3_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i13.GSR = "ENABLED";
    FD1P3AX Out3_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i14.GSR = "ENABLED";
    FD1P3AX Out3_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i15.GSR = "ENABLED";
    FD1P3AX Out3_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i16.GSR = "ENABLED";
    FD1P3AX Out3_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i17.GSR = "ENABLED";
    FD1P3AX Out3_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i18.GSR = "ENABLED";
    FD1P3AX Out3_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i19.GSR = "ENABLED";
    FD1P3AX Out3_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i20.GSR = "ENABLED";
    FD1P3AX Out3_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i21.GSR = "ENABLED";
    FD1P3AX Out3_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i22.GSR = "ENABLED";
    FD1P3AX Out3_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i23.GSR = "ENABLED";
    FD1P3AX Out3_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i24.GSR = "ENABLED";
    FD1P3AX Out3_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i25.GSR = "ENABLED";
    FD1P3AX Out3_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i26.GSR = "ENABLED";
    FD1P3AX Out3_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i27.GSR = "ENABLED";
    FD1P3AX Out3_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_192), 
            .CK(clk_N_875), .Q(Out3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i28.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_220), 
            .CK(clk_N_875), .Q(backOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i1 (.D(backOut3_28__N_1872[1]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i2 (.D(backOut3_28__N_1872[2]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i3 (.D(backOut3_28__N_1872[3]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i4 (.D(backOut3_28__N_1872[4]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i5 (.D(Out2_28__N_1145[5]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i6 (.D(backOut3_28__N_1872[6]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i7 (.D(backOut3_28__N_1872[7]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i8 (.D(backOut3_28__N_1872[8]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i9 (.D(backOut3_28__N_1872[9]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i10 (.D(Out2_28__N_1145[10]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i12 (.D(Out2_28__N_1145[12]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i13 (.D(backOut3_28__N_1872[13]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i14 (.D(backOut3_28__N_1872[14]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i15 (.D(Out2_28__N_1145[15]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i16 (.D(Out2_28__N_1145[16]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i18 (.D(Out2_28__N_1145[18]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i19 (.D(backOut3_28__N_1872[19]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i20 (.D(backOut3_28__N_1872[20]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i21 (.D(Out2_28__N_1145[21]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i22 (.D(backOut3_28__N_1872[22]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i23 (.D(Out0_28__N_1087[23]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i24 (.D(backOut3_28__N_1872[24]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i25 (.D(Out0_28__N_1087[25]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i26 (.D(backOut3_28__N_1872[26]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i28 (.D(Out0_28__N_1087[28]), .SP(clk_N_875_enable_248), 
            .CK(clk_N_875), .Q(backOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i28.GSR = "DISABLED";
    LUT4 mux_189_i9_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[8]), 
         .Z(intgOut0_28__N_1627[8])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i9_3_lut_3_lut.init = 16'hbaba;
    LUT4 mux_189_i7_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[6]), 
         .Z(intgOut0_28__N_1627[6])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i7_3_lut_3_lut.init = 16'hbaba;
    FD1S3AX subOut_i1 (.D(\subOut_24__N_1369[1] ), .CK(clk_N_875), .Q(subOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i1.GSR = "ENABLED";
    FD1S3AX subOut_i2 (.D(\subOut_24__N_1369[2] ), .CK(clk_N_875), .Q(subOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i2.GSR = "ENABLED";
    FD1S3AX subOut_i3 (.D(\subOut_24__N_1369[3] ), .CK(clk_N_875), .Q(subOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i3.GSR = "ENABLED";
    FD1S3AX subOut_i4 (.D(\subOut_24__N_1369[4] ), .CK(clk_N_875), .Q(subOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i4.GSR = "ENABLED";
    FD1S3AX subOut_i5 (.D(\subOut_24__N_1369[5] ), .CK(clk_N_875), .Q(subOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i5.GSR = "ENABLED";
    FD1S3AX subOut_i6 (.D(\subOut_24__N_1369[6] ), .CK(clk_N_875), .Q(subOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i6.GSR = "ENABLED";
    FD1S3AX subOut_i7 (.D(\subOut_24__N_1369[7] ), .CK(clk_N_875), .Q(subOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i7.GSR = "ENABLED";
    FD1S3AX subOut_i8 (.D(\subOut_24__N_1369[8] ), .CK(clk_N_875), .Q(subOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i8.GSR = "ENABLED";
    FD1S3AX subOut_i9 (.D(\subOut_24__N_1369[9] ), .CK(clk_N_875), .Q(subOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i9.GSR = "ENABLED";
    FD1S3AX subOut_i10 (.D(\subOut_24__N_1369[10] ), .CK(clk_N_875), .Q(subOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i10.GSR = "ENABLED";
    FD1S3AX subOut_i11 (.D(\subOut_24__N_1369[11] ), .CK(clk_N_875), .Q(subOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i11.GSR = "ENABLED";
    FD1S3AX subOut_i12 (.D(\subOut_24__N_1369[12] ), .CK(clk_N_875), .Q(subOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i12.GSR = "ENABLED";
    FD1S3AX subOut_i13 (.D(\subOut_24__N_1369[13] ), .CK(clk_N_875), .Q(subOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i13.GSR = "ENABLED";
    FD1S3AX subOut_i14 (.D(\subOut_24__N_1369[14] ), .CK(clk_N_875), .Q(subOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i14.GSR = "ENABLED";
    FD1S3AX subOut_i15 (.D(\subOut_24__N_1369[15] ), .CK(clk_N_875), .Q(subOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i15.GSR = "ENABLED";
    FD1S3AX subOut_i16 (.D(\subOut_24__N_1369[16] ), .CK(clk_N_875), .Q(subOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i16.GSR = "ENABLED";
    FD1S3AX subOut_i17 (.D(\subOut_24__N_1369[17] ), .CK(clk_N_875), .Q(subOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i17.GSR = "ENABLED";
    FD1S3AX subOut_i18 (.D(\subOut_24__N_1369[18] ), .CK(clk_N_875), .Q(subOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i18.GSR = "ENABLED";
    FD1S3AX subOut_i19 (.D(\subOut_24__N_1369[19] ), .CK(clk_N_875), .Q(subOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i19.GSR = "ENABLED";
    FD1S3AX subOut_i20 (.D(\subOut_24__N_1369[20] ), .CK(clk_N_875), .Q(subOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i20.GSR = "ENABLED";
    FD1S3AX subOut_i21 (.D(\subOut_24__N_1369[21] ), .CK(clk_N_875), .Q(subOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i21.GSR = "ENABLED";
    FD1S3AX subOut_i23 (.D(\subOut_24__N_1369[24] ), .CK(clk_N_875), .Q(subOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i23.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_68 (.A(n16481), .B(n16131), .C(n21677), .D(n22440), 
         .Z(clk_N_875_enable_389)) /* synthesis lut_function=((B (C (D))+!B (C+!(D)))+!A) */ ;
    defparam i1_4_lut_adj_68.init = 16'hf577;
    LUT4 i13137_2_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[5]), .Z(intgOut0_28__N_1627[5])) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i13137_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_69 (.A(n3612), .B(n35_adj_2342), .C(n40_adj_2343), 
         .D(n36_adj_2344), .Z(n4_adj_2341)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_69.init = 16'haaa8;
    LUT4 i14_4_lut_adj_70 (.A(speed_set_m1[13]), .B(speed_set_m1[1]), .C(speed_set_m1[12]), 
         .D(speed_set_m1[2]), .Z(n35_adj_2342)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_70.init = 16'hfffe;
    LUT4 i19_4_lut_adj_71 (.A(speed_set_m1[15]), .B(n38_adj_2345), .C(n32_adj_2346), 
         .D(speed_set_m1[10]), .Z(n40_adj_2343)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_71.init = 16'hfffe;
    LUT4 i15_4_lut_adj_72 (.A(speed_set_m1[0]), .B(speed_set_m1[7]), .C(speed_set_m1[17]), 
         .D(speed_set_m1[11]), .Z(n36_adj_2344)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_72.init = 16'hfffe;
    LUT4 i17_4_lut_adj_73 (.A(speed_set_m1[8]), .B(n34_adj_2347), .C(n24_adj_2348), 
         .D(speed_set_m1[16]), .Z(n38_adj_2345)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_73.init = 16'hfffe;
    LUT4 i11_3_lut_adj_74 (.A(speed_set_m1[6]), .B(speed_set_m1[3]), .C(speed_set_m1[14]), 
         .Z(n32_adj_2346)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_74.init = 16'hfefe;
    CCU2D add_15370_5 (.A0(addOut[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18756), .COUT(n18757));
    defparam add_15370_5.INIT0 = 16'hf555;
    defparam add_15370_5.INIT1 = 16'h0aaa;
    defparam add_15370_5.INJECT1_0 = "NO";
    defparam add_15370_5.INJECT1_1 = "NO";
    CCU2D add_15370_3 (.A0(addOut[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18755), .COUT(n18756));
    defparam add_15370_3.INIT0 = 16'hf555;
    defparam add_15370_3.INIT1 = 16'hf555;
    defparam add_15370_3.INJECT1_0 = "NO";
    defparam add_15370_3.INJECT1_1 = "NO";
    LUT4 i13_4_lut_adj_75 (.A(speed_set_m1[20]), .B(speed_set_m1[19]), .C(speed_set_m1[9]), 
         .D(speed_set_m1[4]), .Z(n34_adj_2347)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_75.init = 16'hfffe;
    CCU2D add_15370_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[0]), .B1(addOut[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18755));
    defparam add_15370_1.INIT0 = 16'hF000;
    defparam add_15370_1.INIT1 = 16'ha666;
    defparam add_15370_1.INJECT1_0 = "NO";
    defparam add_15370_1.INJECT1_1 = "NO";
    CCU2D add_15378_9 (.A0(speed_set_m1[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18642), .COUT(n18643));
    defparam add_15378_9.INIT0 = 16'hf555;
    defparam add_15378_9.INIT1 = 16'h0aaa;
    defparam add_15378_9.INJECT1_0 = "NO";
    defparam add_15378_9.INJECT1_1 = "NO";
    LUT4 i3_2_lut_adj_76 (.A(speed_set_m1[18]), .B(speed_set_m1[5]), .Z(n24_adj_2348)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_76.init = 16'heeee;
    LUT4 i1_4_lut_4_lut_adj_77 (.A(n21630), .B(n16073), .C(n21636), .D(n21631), 
         .Z(n19942)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam i1_4_lut_4_lut_adj_77.init = 16'h5400;
    LUT4 mux_135_i24_4_lut (.A(backOut2[23]), .B(backOut3[23]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i24_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_78 (.A(ss[2]), .B(n19907), .C(n22440), .D(n4_adj_2349), 
         .Z(clk_N_875_enable_72)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_78.init = 16'hc8c0;
    LUT4 i1_3_lut_adj_79 (.A(ss[0]), .B(ss[3]), .C(ss[1]), .Z(n4_adj_2349)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_3_lut_adj_79.init = 16'h0202;
    LUT4 mux_135_i25_4_lut (.A(backOut2[24]), .B(backOut3[24]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i25_4_lut.init = 16'h0aca;
    LUT4 i2_3_lut_4_lut (.A(n21633), .B(n21632), .C(subIn1_24__N_1342), 
         .D(n21637), .Z(n11474)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0800;
    LUT4 mux_135_i2_4_lut (.A(backOut2[1]), .B(backOut3[1]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i2_4_lut.init = 16'h0aca;
    LUT4 i7_4_lut (.A(Out3[3]), .B(n14_adj_2350), .C(n10), .D(Out3[4]), 
         .Z(n18960)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut (.A(Out3[11]), .B(Out3[7]), .C(Out3[2]), .D(Out3[10]), 
         .Z(n14_adj_2350)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(Out3[9]), .B(Out3[1]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i4_4_lut (.A(Out3[5]), .B(Out3[6]), .C(Out3[0]), .D(n6_adj_2351), 
         .Z(n18961)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_80 (.A(Out3[8]), .B(Out3[12]), .Z(n6_adj_2351)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i1_2_lut_adj_80.init = 16'heeee;
    LUT4 mux_135_i26_4_lut (.A(backOut2[25]), .B(backOut3[25]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i26_4_lut.init = 16'h0aca;
    LUT4 mux_135_i3_4_lut (.A(backOut2[2]), .B(backOut3[2]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i3_4_lut.init = 16'h0aca;
    LUT4 mux_135_i27_4_lut (.A(backOut2[26]), .B(backOut3[26]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i27_4_lut.init = 16'h0aca;
    LUT4 mux_135_i4_4_lut (.A(backOut2[3]), .B(backOut3[3]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i4_4_lut.init = 16'h0aca;
    LUT4 mux_135_i28_4_lut (.A(backOut2[27]), .B(backOut3[27]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i28_4_lut.init = 16'h0aca;
    LUT4 mux_135_i5_4_lut (.A(backOut2[4]), .B(backOut3[4]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i5_4_lut.init = 16'h0aca;
    LUT4 mux_135_i29_4_lut (.A(backOut2[28]), .B(backOut3[28]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i29_4_lut.init = 16'h0aca;
    LUT4 mux_135_i6_4_lut (.A(backOut2[5]), .B(backOut3[5]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i6_4_lut.init = 16'h0aca;
    LUT4 mux_135_i7_4_lut (.A(backOut2[6]), .B(backOut3[6]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i7_4_lut.init = 16'h0aca;
    LUT4 i13138_2_lut (.A(addOut[0]), .B(n22440), .Z(Out3_28__N_1174[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13138_2_lut.init = 16'h2222;
    LUT4 mux_135_i8_4_lut (.A(backOut2[7]), .B(backOut3[7]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i8_4_lut.init = 16'h0aca;
    LUT4 mux_135_i1_4_lut (.A(backOut2[0]), .B(backOut3[0]), .C(n21659), 
         .D(n9_adj_2331), .Z(n555[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i1_4_lut.init = 16'h0aca;
    LUT4 i7_4_lut_adj_81 (.A(Out0[3]), .B(n14_adj_2352), .C(n10_adj_2353), 
         .D(Out0[4]), .Z(n18945)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i7_4_lut_adj_81.init = 16'hfffe;
    LUT4 i6_4_lut_adj_82 (.A(Out0[11]), .B(Out0[7]), .C(Out0[2]), .D(Out0[10]), 
         .Z(n14_adj_2352)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i6_4_lut_adj_82.init = 16'hfffe;
    LUT4 i2_2_lut_adj_83 (.A(Out0[9]), .B(Out0[1]), .Z(n10_adj_2353)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i2_2_lut_adj_83.init = 16'heeee;
    LUT4 i4_4_lut_adj_84 (.A(Out0[5]), .B(Out0[6]), .C(Out0[0]), .D(n6_adj_2354), 
         .Z(n18946)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i4_4_lut_adj_84.init = 16'hfffe;
    LUT4 i1_2_lut_adj_85 (.A(Out0[8]), .B(Out0[12]), .Z(n6_adj_2354)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i1_2_lut_adj_85.init = 16'heeee;
    LUT4 i7_4_lut_adj_86 (.A(Out1[3]), .B(n14_adj_2355), .C(n10_adj_2356), 
         .D(Out1[4]), .Z(n18920)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i7_4_lut_adj_86.init = 16'hfffe;
    LUT4 i6_4_lut_adj_87 (.A(Out1[11]), .B(Out1[7]), .C(Out1[2]), .D(Out1[10]), 
         .Z(n14_adj_2355)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i6_4_lut_adj_87.init = 16'hfffe;
    LUT4 i2_2_lut_adj_88 (.A(Out1[9]), .B(Out1[1]), .Z(n10_adj_2356)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i2_2_lut_adj_88.init = 16'heeee;
    LUT4 i4_4_lut_adj_89 (.A(Out1[5]), .B(Out1[6]), .C(Out1[0]), .D(n6_adj_2357), 
         .Z(n18921)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i4_4_lut_adj_89.init = 16'hfffe;
    LUT4 i1_2_lut_adj_90 (.A(Out1[8]), .B(Out1[12]), .Z(n6_adj_2357)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i1_2_lut_adj_90.init = 16'heeee;
    LUT4 i17460_4_lut (.A(ss[3]), .B(ss[0]), .C(ss[2]), .D(n22440), 
         .Z(n16283)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+((D)+!C))) */ ;
    defparam i17460_4_lut.init = 16'hffed;
    LUT4 i11751_4_lut (.A(clk_N_875_enable_391), .B(n1294[15]), .C(n9), 
         .D(n18943), .Z(n14336)) /* synthesis lut_function=(A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11751_4_lut.init = 16'haa2a;
    LUT4 i1_2_lut_rep_345_4_lut (.A(n22440), .B(n21697), .C(ss[3]), .D(ss[0]), 
         .Z(n21658)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(164[13] 176[6])
    defparam i1_2_lut_rep_345_4_lut.init = 16'h1400;
    LUT4 i5_4_lut (.A(n9_adj_2358), .B(n1294[10]), .C(n8), .D(n1294[11]), 
         .Z(n9)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i3_2_lut_adj_91 (.A(n1294[14]), .B(n1294[13]), .Z(n9_adj_2358)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_91.init = 16'h8888;
    LUT4 i2_4_lut_adj_92 (.A(n1294[9]), .B(n1294[12]), .C(n10_adj_2359), 
         .D(n1294[7]), .Z(n8)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_92.init = 16'hccc8;
    LUT4 i1_4_lut_adj_93 (.A(ss[3]), .B(n19907), .C(n22440), .D(n21676), 
         .Z(clk_N_875_enable_44)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_93.init = 16'hc4c0;
    LUT4 i4_4_lut_adj_94 (.A(n1294[6]), .B(n8_adj_2360), .C(n1294[4]), 
         .D(n4_adj_2361), .Z(n10_adj_2359)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_94.init = 16'hfeee;
    LUT4 i2_2_lut_adj_95 (.A(n1294[5]), .B(n1294[8]), .Z(n8_adj_2360)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_95.init = 16'heeee;
    LUT4 i1_4_lut_adj_96 (.A(n1294[3]), .B(n1294[2]), .C(n1294[1]), .D(n1294[0]), 
         .Z(n4_adj_2361)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_96.init = 16'haaa8;
    CCU2D add_15378_7 (.A0(speed_set_m1[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18641), .COUT(n18642));
    defparam add_15378_7.INIT0 = 16'h0aaa;
    defparam add_15378_7.INIT1 = 16'hf555;
    defparam add_15378_7.INJECT1_0 = "NO";
    defparam add_15378_7.INJECT1_1 = "NO";
    CCU2D add_15378_5 (.A0(speed_set_m1[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18640), .COUT(n18641));
    defparam add_15378_5.INIT0 = 16'h0aaa;
    defparam add_15378_5.INIT1 = 16'h0aaa;
    defparam add_15378_5.INJECT1_0 = "NO";
    defparam add_15378_5.INJECT1_1 = "NO";
    CCU2D add_15378_3 (.A0(speed_set_m1[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18639), .COUT(n18640));
    defparam add_15378_3.INIT0 = 16'hf555;
    defparam add_15378_3.INIT1 = 16'hf555;
    defparam add_15378_3.INJECT1_0 = "NO";
    defparam add_15378_3.INJECT1_1 = "NO";
    CCU2D add_15378_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[4]), .B1(speed_set_m1[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18639));
    defparam add_15378_1.INIT0 = 16'hF000;
    defparam add_15378_1.INIT1 = 16'ha666;
    defparam add_15378_1.INJECT1_0 = "NO";
    defparam add_15378_1.INJECT1_1 = "NO";
    CCU2D add_15379_21 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18638), .S1(n49));
    defparam add_15379_21.INIT0 = 16'h5555;
    defparam add_15379_21.INIT1 = 16'h0000;
    defparam add_15379_21.INJECT1_0 = "NO";
    defparam add_15379_21.INJECT1_1 = "NO";
    CCU2D add_15379_19 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18637), .COUT(n18638));
    defparam add_15379_19.INIT0 = 16'hf555;
    defparam add_15379_19.INIT1 = 16'hf555;
    defparam add_15379_19.INJECT1_0 = "NO";
    defparam add_15379_19.INJECT1_1 = "NO";
    CCU2D add_15379_17 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18636), .COUT(n18637));
    defparam add_15379_17.INIT0 = 16'hf555;
    defparam add_15379_17.INIT1 = 16'hf555;
    defparam add_15379_17.INJECT1_0 = "NO";
    defparam add_15379_17.INJECT1_1 = "NO";
    CCU2D add_15379_15 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18635), .COUT(n18636));
    defparam add_15379_15.INIT0 = 16'hf555;
    defparam add_15379_15.INIT1 = 16'hf555;
    defparam add_15379_15.INJECT1_0 = "NO";
    defparam add_15379_15.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_97 (.A(ss[0]), .B(n21694), .C(ss[3]), .D(n22440), 
         .Z(n19947)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_3_lut_4_lut_adj_97.init = 16'h0080;
    CCU2D add_223_11 (.A0(Out3[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18449), 
          .COUT(n18450), .S0(n1357[9]), .S1(n1357[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_11.INIT0 = 16'h5aaa;
    defparam add_223_11.INIT1 = 16'h5aaa;
    defparam add_223_11.INJECT1_0 = "NO";
    defparam add_223_11.INJECT1_1 = "NO";
    CCU2D add_15379_13 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18634), .COUT(n18635));
    defparam add_15379_13.INIT0 = 16'hf555;
    defparam add_15379_13.INIT1 = 16'hf555;
    defparam add_15379_13.INJECT1_0 = "NO";
    defparam add_15379_13.INJECT1_1 = "NO";
    CCU2D add_15379_11 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18633), .COUT(n18634));
    defparam add_15379_11.INIT0 = 16'hf555;
    defparam add_15379_11.INIT1 = 16'hf555;
    defparam add_15379_11.INJECT1_0 = "NO";
    defparam add_15379_11.INJECT1_1 = "NO";
    CCU2D add_211_15 (.A0(Out0[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18427), 
          .COUT(n18428), .S0(n1294[13]), .S1(n1294[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_15.INIT0 = 16'h5aaa;
    defparam add_211_15.INIT1 = 16'h5aaa;
    defparam add_211_15.INJECT1_0 = "NO";
    defparam add_211_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_98 (.A(n21698), .B(n21697), .C(n22435), 
         .D(n22440), .Z(n19907)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut_4_lut_adj_98.init = 16'he0f0;
    CCU2D add_211_13 (.A0(Out0[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18426), 
          .COUT(n18427), .S0(n1294[11]), .S1(n1294[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_13.INIT0 = 16'h5aaa;
    defparam add_211_13.INIT1 = 16'h5aaa;
    defparam add_211_13.INJECT1_0 = "NO";
    defparam add_211_13.INJECT1_1 = "NO";
    LUT4 i11671_3_lut_4_lut (.A(ss[2]), .B(n21698), .C(n19967), .D(clk_N_875_enable_389), 
         .Z(n14237)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11671_3_lut_4_lut.init = 16'hfd00;
    CCU2D add_15379_9 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18632), .COUT(n18633));
    defparam add_15379_9.INIT0 = 16'hf555;
    defparam add_15379_9.INIT1 = 16'hf555;
    defparam add_15379_9.INJECT1_0 = "NO";
    defparam add_15379_9.INJECT1_1 = "NO";
    LUT4 mux_138_i15_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[14]), 
         .D(intgOut2[14]), .Z(n645[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 i11699_3_lut_4_lut (.A(ss[2]), .B(n21698), .C(n19964), .D(clk_N_875_enable_392), 
         .Z(n14265)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11699_3_lut_4_lut.init = 16'hfd00;
    CCU2D add_15379_7 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18631), .COUT(n18632));
    defparam add_15379_7.INIT0 = 16'hf555;
    defparam add_15379_7.INIT1 = 16'hf555;
    defparam add_15379_7.INJECT1_0 = "NO";
    defparam add_15379_7.INJECT1_1 = "NO";
    CCU2D add_15379_5 (.A0(speed_set_m3[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18630), .COUT(n18631));
    defparam add_15379_5.INIT0 = 16'hf555;
    defparam add_15379_5.INIT1 = 16'hf555;
    defparam add_15379_5.INJECT1_0 = "NO";
    defparam add_15379_5.INJECT1_1 = "NO";
    CCU2D add_15379_3 (.A0(speed_set_m3[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18629), .COUT(n18630));
    defparam add_15379_3.INIT0 = 16'hf555;
    defparam add_15379_3.INIT1 = 16'hf555;
    defparam add_15379_3.INJECT1_0 = "NO";
    defparam add_15379_3.INJECT1_1 = "NO";
    CCU2D add_15388_21 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18736), .S1(n56));
    defparam add_15388_21.INIT0 = 16'h5555;
    defparam add_15388_21.INIT1 = 16'h0000;
    defparam add_15388_21.INJECT1_0 = "NO";
    defparam add_15388_21.INJECT1_1 = "NO";
    CCU2D add_15379_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[0]), .B1(speed_set_m3[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18629));
    defparam add_15379_1.INIT0 = 16'hF000;
    defparam add_15379_1.INIT1 = 16'ha666;
    defparam add_15379_1.INJECT1_0 = "NO";
    defparam add_15379_1.INJECT1_1 = "NO";
    CCU2D add_15388_19 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18735), .COUT(n18736));
    defparam add_15388_19.INIT0 = 16'hf555;
    defparam add_15388_19.INIT1 = 16'hf555;
    defparam add_15388_19.INJECT1_0 = "NO";
    defparam add_15388_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_420 (.A(n22440), .B(n22433), .C(ss[3]), .Z(n22424)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam i1_2_lut_rep_420.init = 16'hfbfb;
    LUT4 i11760_4_lut (.A(clk_N_875_enable_391), .B(n18943), .C(n30), 
         .D(n1315[15]), .Z(n14345)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11760_4_lut.init = 16'h8aaa;
    LUT4 i5_4_lut_adj_99 (.A(n9_adj_2362), .B(n7), .C(n1315[10]), .D(n1315[13]), 
         .Z(n30)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_99.init = 16'h8000;
    LUT4 i3_2_lut_adj_100 (.A(n1315[14]), .B(n1315[12]), .Z(n9_adj_2362)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_100.init = 16'h8888;
    LUT4 i1_4_lut_adj_101 (.A(n1315[11]), .B(n1315[9]), .C(n10_adj_2363), 
         .D(n1315[7]), .Z(n7)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_101.init = 16'haaa8;
    CCU2D add_15388_17 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18734), .COUT(n18735));
    defparam add_15388_17.INIT0 = 16'hf555;
    defparam add_15388_17.INIT1 = 16'hf555;
    defparam add_15388_17.INJECT1_0 = "NO";
    defparam add_15388_17.INJECT1_1 = "NO";
    LUT4 i4_4_lut_adj_102 (.A(n1315[6]), .B(n8_adj_2364), .C(n1315[4]), 
         .D(n4_adj_2365), .Z(n10_adj_2363)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_102.init = 16'hfeee;
    LUT4 i2_2_lut_adj_103 (.A(n1315[5]), .B(n1315[8]), .Z(n8_adj_2364)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_103.init = 16'heeee;
    CCU2D add_15380_21 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18628), .S1(n42));
    defparam add_15380_21.INIT0 = 16'h5555;
    defparam add_15380_21.INIT1 = 16'h0000;
    defparam add_15380_21.INJECT1_0 = "NO";
    defparam add_15380_21.INJECT1_1 = "NO";
    CCU2D add_15380_19 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18627), .COUT(n18628));
    defparam add_15380_19.INIT0 = 16'hf555;
    defparam add_15380_19.INIT1 = 16'hf555;
    defparam add_15380_19.INJECT1_0 = "NO";
    defparam add_15380_19.INJECT1_1 = "NO";
    CCU2D add_15380_17 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18626), .COUT(n18627));
    defparam add_15380_17.INIT0 = 16'hf555;
    defparam add_15380_17.INIT1 = 16'hf555;
    defparam add_15380_17.INJECT1_0 = "NO";
    defparam add_15380_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_104 (.A(n1315[3]), .B(n1315[2]), .C(n1315[1]), .D(n1315[0]), 
         .Z(n4_adj_2365)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_104.init = 16'haaa8;
    LUT4 i13254_2_lut (.A(addOut[8]), .B(n22440), .Z(backOut3_28__N_1872[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13254_2_lut.init = 16'h2222;
    LUT4 i13253_2_lut (.A(addOut[7]), .B(n22440), .Z(backOut3_28__N_1872[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13253_2_lut.init = 16'h2222;
    LUT4 i13252_2_lut (.A(addOut[6]), .B(n22440), .Z(backOut3_28__N_1872[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13252_2_lut.init = 16'h2222;
    LUT4 i13459_2_lut (.A(addOut[5]), .B(n22440), .Z(Out2_28__N_1145[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13459_2_lut.init = 16'h2222;
    LUT4 i13250_2_lut (.A(addOut[4]), .B(n22440), .Z(backOut3_28__N_1872[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13250_2_lut.init = 16'h2222;
    LUT4 i13249_2_lut (.A(addOut[3]), .B(n22440), .Z(backOut3_28__N_1872[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13249_2_lut.init = 16'h2222;
    LUT4 i13248_2_lut (.A(addOut[2]), .B(n22440), .Z(backOut3_28__N_1872[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13248_2_lut.init = 16'h2222;
    LUT4 i13247_2_lut (.A(addOut[1]), .B(n22440), .Z(backOut3_28__N_1872[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13247_2_lut.init = 16'h2222;
    LUT4 i11747_3_lut_4_lut (.A(ss[2]), .B(n21728), .C(n19964), .D(clk_N_875_enable_309), 
         .Z(n14313)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11747_3_lut_4_lut.init = 16'hfe00;
    LUT4 i11723_3_lut_4_lut (.A(ss[2]), .B(n21728), .C(n19967), .D(clk_N_875_enable_333), 
         .Z(n14289)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11723_3_lut_4_lut.init = 16'hfe00;
    LUT4 i17532_2_lut_3_lut_4_lut (.A(n21729), .B(n22419), .C(n22423), 
         .D(ss[2]), .Z(n20659)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i17532_2_lut_3_lut_4_lut.init = 16'hf0f4;
    CCU2D add_15380_15 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18625), .COUT(n18626));
    defparam add_15380_15.INIT0 = 16'hf555;
    defparam add_15380_15.INIT1 = 16'hf555;
    defparam add_15380_15.INJECT1_0 = "NO";
    defparam add_15380_15.INJECT1_1 = "NO";
    CCU2D add_15380_13 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18624), .COUT(n18625));
    defparam add_15380_13.INIT0 = 16'hf555;
    defparam add_15380_13.INIT1 = 16'hf555;
    defparam add_15380_13.INJECT1_0 = "NO";
    defparam add_15380_13.INJECT1_1 = "NO";
    CCU2D add_15388_15 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18733), .COUT(n18734));
    defparam add_15388_15.INIT0 = 16'hf555;
    defparam add_15388_15.INIT1 = 16'hf555;
    defparam add_15388_15.INJECT1_0 = "NO";
    defparam add_15388_15.INJECT1_1 = "NO";
    CCU2D add_15388_13 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18732), .COUT(n18733));
    defparam add_15388_13.INIT0 = 16'hf555;
    defparam add_15388_13.INIT1 = 16'hf555;
    defparam add_15388_13.INJECT1_0 = "NO";
    defparam add_15388_13.INJECT1_1 = "NO";
    CCU2D add_15380_11 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18623), .COUT(n18624));
    defparam add_15380_11.INIT0 = 16'hf555;
    defparam add_15380_11.INIT1 = 16'hf555;
    defparam add_15380_11.INJECT1_0 = "NO";
    defparam add_15380_11.INJECT1_1 = "NO";
    CCU2D add_223_9 (.A0(Out3[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18448), 
          .COUT(n18449), .S0(n1357[7]), .S1(n1357[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_9.INIT0 = 16'h5aaa;
    defparam add_223_9.INIT1 = 16'h5aaa;
    defparam add_223_9.INJECT1_0 = "NO";
    defparam add_223_9.INJECT1_1 = "NO";
    CCU2D add_15380_9 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18622), .COUT(n18623));
    defparam add_15380_9.INIT0 = 16'hf555;
    defparam add_15380_9.INIT1 = 16'hf555;
    defparam add_15380_9.INJECT1_0 = "NO";
    defparam add_15380_9.INJECT1_1 = "NO";
    CCU2D add_15388_11 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18731), .COUT(n18732));
    defparam add_15388_11.INIT0 = 16'hf555;
    defparam add_15388_11.INIT1 = 16'hf555;
    defparam add_15388_11.INJECT1_0 = "NO";
    defparam add_15388_11.INJECT1_1 = "NO";
    CCU2D add_15388_9 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18730), .COUT(n18731));
    defparam add_15388_9.INIT0 = 16'hf555;
    defparam add_15388_9.INIT1 = 16'hf555;
    defparam add_15388_9.INJECT1_0 = "NO";
    defparam add_15388_9.INJECT1_1 = "NO";
    CCU2D add_15388_7 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18729), .COUT(n18730));
    defparam add_15388_7.INIT0 = 16'hf555;
    defparam add_15388_7.INIT1 = 16'hf555;
    defparam add_15388_7.INJECT1_0 = "NO";
    defparam add_15388_7.INJECT1_1 = "NO";
    CCU2D add_15388_5 (.A0(speed_set_m4[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18728), .COUT(n18729));
    defparam add_15388_5.INIT0 = 16'hf555;
    defparam add_15388_5.INIT1 = 16'hf555;
    defparam add_15388_5.INJECT1_0 = "NO";
    defparam add_15388_5.INJECT1_1 = "NO";
    CCU2D add_15388_3 (.A0(speed_set_m4[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18727), .COUT(n18728));
    defparam add_15388_3.INIT0 = 16'hf555;
    defparam add_15388_3.INIT1 = 16'hf555;
    defparam add_15388_3.INJECT1_0 = "NO";
    defparam add_15388_3.INJECT1_1 = "NO";
    CCU2D add_15380_7 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18621), .COUT(n18622));
    defparam add_15380_7.INIT0 = 16'hf555;
    defparam add_15380_7.INIT1 = 16'hf555;
    defparam add_15380_7.INJECT1_0 = "NO";
    defparam add_15380_7.INJECT1_1 = "NO";
    CCU2D add_15388_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[0]), .B1(speed_set_m4[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18727));
    defparam add_15388_1.INIT0 = 16'hF000;
    defparam add_15388_1.INIT1 = 16'ha666;
    defparam add_15388_1.INJECT1_0 = "NO";
    defparam add_15388_1.INJECT1_1 = "NO";
    CCU2D add_223_7 (.A0(Out3[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18447), 
          .COUT(n18448), .S0(n1357[5]), .S1(n1357[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_7.INIT0 = 16'h5aaa;
    defparam add_223_7.INIT1 = 16'h5aaa;
    defparam add_223_7.INJECT1_0 = "NO";
    defparam add_223_7.INJECT1_1 = "NO";
    PFUMX i17827 (.BLUT(n22426), .ALUT(n22427), .C0(ss[0]), .Z(n21648));
    CCU2D add_15371_24 (.A0(addOut[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18726), 
          .S1(n1065));
    defparam add_15371_24.INIT0 = 16'hf555;
    defparam add_15371_24.INIT1 = 16'h0000;
    defparam add_15371_24.INJECT1_0 = "NO";
    defparam add_15371_24.INJECT1_1 = "NO";
    CCU2D add_223_5 (.A0(Out3[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18446), 
          .COUT(n18447), .S0(n1357[3]), .S1(n1357[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_5.INIT0 = 16'h5aaa;
    defparam add_223_5.INIT1 = 16'h5aaa;
    defparam add_223_5.INJECT1_0 = "NO";
    defparam add_223_5.INJECT1_1 = "NO";
    LUT4 i13580_2_lut_rep_320 (.A(n15564), .B(n49), .Z(n21633)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13580_2_lut_rep_320.init = 16'heeee;
    CCU2D add_223_3 (.A0(Out3[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18445), 
          .COUT(n18446), .S0(n1357[1]), .S1(n1357[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_3.INIT0 = 16'h5aaa;
    defparam add_223_3.INIT1 = 16'h5aaa;
    defparam add_223_3.INJECT1_0 = "NO";
    defparam add_223_3.INJECT1_1 = "NO";
    CCU2D add_211_11 (.A0(Out0[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18425), 
          .COUT(n18426), .S0(n1294[9]), .S1(n1294[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_11.INIT0 = 16'h5aaa;
    defparam add_211_11.INIT1 = 16'h5aaa;
    defparam add_211_11.INJECT1_0 = "NO";
    defparam add_211_11.INJECT1_1 = "NO";
    CCU2D add_15380_5 (.A0(speed_set_m2[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18620), .COUT(n18621));
    defparam add_15380_5.INIT0 = 16'hf555;
    defparam add_15380_5.INIT1 = 16'hf555;
    defparam add_15380_5.INJECT1_0 = "NO";
    defparam add_15380_5.INJECT1_1 = "NO";
    CCU2D add_15380_3 (.A0(speed_set_m2[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18619), .COUT(n18620));
    defparam add_15380_3.INIT0 = 16'hf555;
    defparam add_15380_3.INIT1 = 16'hf555;
    defparam add_15380_3.INJECT1_0 = "NO";
    defparam add_15380_3.INJECT1_1 = "NO";
    CCU2D add_15371_22 (.A0(addOut[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18725), .COUT(n18726));
    defparam add_15371_22.INIT0 = 16'h5555;
    defparam add_15371_22.INIT1 = 16'h5555;
    defparam add_15371_22.INJECT1_0 = "NO";
    defparam add_15371_22.INJECT1_1 = "NO";
    CCU2D add_15380_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[0]), .B1(speed_set_m2[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18619));
    defparam add_15380_1.INIT0 = 16'hF000;
    defparam add_15380_1.INIT1 = 16'ha666;
    defparam add_15380_1.INJECT1_0 = "NO";
    defparam add_15380_1.INJECT1_1 = "NO";
    CCU2D add_15381_21 (.A0(speed_set_m1[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18618), .S1(n35));
    defparam add_15381_21.INIT0 = 16'h5555;
    defparam add_15381_21.INIT1 = 16'h0000;
    defparam add_15381_21.INJECT1_0 = "NO";
    defparam add_15381_21.INJECT1_1 = "NO";
    CCU2D add_15381_19 (.A0(speed_set_m1[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18617), .COUT(n18618));
    defparam add_15381_19.INIT0 = 16'hf555;
    defparam add_15381_19.INIT1 = 16'hf555;
    defparam add_15381_19.INJECT1_0 = "NO";
    defparam add_15381_19.INJECT1_1 = "NO";
    CCU2D add_15371_20 (.A0(addOut[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18724), .COUT(n18725));
    defparam add_15371_20.INIT0 = 16'h5555;
    defparam add_15371_20.INIT1 = 16'h5555;
    defparam add_15371_20.INJECT1_0 = "NO";
    defparam add_15371_20.INJECT1_1 = "NO";
    CCU2D add_15371_18 (.A0(addOut[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18723), .COUT(n18724));
    defparam add_15371_18.INIT0 = 16'h5555;
    defparam add_15371_18.INIT1 = 16'h5555;
    defparam add_15371_18.INJECT1_0 = "NO";
    defparam add_15371_18.INJECT1_1 = "NO";
    CCU2D add_15371_16 (.A0(addOut[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18722), .COUT(n18723));
    defparam add_15371_16.INIT0 = 16'h5aaa;
    defparam add_15371_16.INIT1 = 16'h5555;
    defparam add_15371_16.INJECT1_0 = "NO";
    defparam add_15371_16.INJECT1_1 = "NO";
    CCU2D add_15381_17 (.A0(speed_set_m1[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18616), .COUT(n18617));
    defparam add_15381_17.INIT0 = 16'hf555;
    defparam add_15381_17.INIT1 = 16'hf555;
    defparam add_15381_17.INJECT1_0 = "NO";
    defparam add_15381_17.INJECT1_1 = "NO";
    CCU2D add_15381_15 (.A0(speed_set_m1[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18615), .COUT(n18616));
    defparam add_15381_15.INIT0 = 16'hf555;
    defparam add_15381_15.INIT1 = 16'hf555;
    defparam add_15381_15.INJECT1_0 = "NO";
    defparam add_15381_15.INJECT1_1 = "NO";
    CCU2D add_15381_13 (.A0(speed_set_m1[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18614), .COUT(n18615));
    defparam add_15381_13.INIT0 = 16'hf555;
    defparam add_15381_13.INIT1 = 16'hf555;
    defparam add_15381_13.INJECT1_0 = "NO";
    defparam add_15381_13.INJECT1_1 = "NO";
    CCU2D add_15381_11 (.A0(speed_set_m1[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18613), .COUT(n18614));
    defparam add_15381_11.INIT0 = 16'hf555;
    defparam add_15381_11.INIT1 = 16'hf555;
    defparam add_15381_11.INJECT1_0 = "NO";
    defparam add_15381_11.INJECT1_1 = "NO";
    CCU2D add_15371_14 (.A0(addOut[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18721), .COUT(n18722));
    defparam add_15371_14.INIT0 = 16'h5aaa;
    defparam add_15371_14.INIT1 = 16'h5555;
    defparam add_15371_14.INJECT1_0 = "NO";
    defparam add_15371_14.INJECT1_1 = "NO";
    CCU2D add_15371_12 (.A0(addOut[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18720), .COUT(n18721));
    defparam add_15371_12.INIT0 = 16'h5555;
    defparam add_15371_12.INIT1 = 16'h5aaa;
    defparam add_15371_12.INJECT1_0 = "NO";
    defparam add_15371_12.INJECT1_1 = "NO";
    CCU2D add_15381_9 (.A0(speed_set_m1[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18612), .COUT(n18613));
    defparam add_15381_9.INIT0 = 16'hf555;
    defparam add_15381_9.INIT1 = 16'hf555;
    defparam add_15381_9.INJECT1_0 = "NO";
    defparam add_15381_9.INJECT1_1 = "NO";
    CCU2D add_15381_7 (.A0(speed_set_m1[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18611), .COUT(n18612));
    defparam add_15381_7.INIT0 = 16'hf555;
    defparam add_15381_7.INIT1 = 16'hf555;
    defparam add_15381_7.INJECT1_0 = "NO";
    defparam add_15381_7.INJECT1_1 = "NO";
    CCU2D add_15381_5 (.A0(speed_set_m1[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18610), .COUT(n18611));
    defparam add_15381_5.INIT0 = 16'hf555;
    defparam add_15381_5.INIT1 = 16'hf555;
    defparam add_15381_5.INJECT1_0 = "NO";
    defparam add_15381_5.INJECT1_1 = "NO";
    CCU2D add_15381_3 (.A0(speed_set_m1[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18609), .COUT(n18610));
    defparam add_15381_3.INIT0 = 16'hf555;
    defparam add_15381_3.INIT1 = 16'hf555;
    defparam add_15381_3.INJECT1_0 = "NO";
    defparam add_15381_3.INJECT1_1 = "NO";
    CCU2D add_15371_10 (.A0(addOut[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18719), .COUT(n18720));
    defparam add_15371_10.INIT0 = 16'h5aaa;
    defparam add_15371_10.INIT1 = 16'h5aaa;
    defparam add_15371_10.INJECT1_0 = "NO";
    defparam add_15371_10.INJECT1_1 = "NO";
    CCU2D add_15371_8 (.A0(addOut[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18718), .COUT(n18719));
    defparam add_15371_8.INIT0 = 16'h5555;
    defparam add_15371_8.INIT1 = 16'h5aaa;
    defparam add_15371_8.INJECT1_0 = "NO";
    defparam add_15371_8.INJECT1_1 = "NO";
    CCU2D add_223_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[13]), .B1(n18960), .C1(n18961), .D1(Out3[28]), .COUT(n18445), 
          .S1(n1357[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_1.INIT0 = 16'hF000;
    defparam add_223_1.INIT1 = 16'h56aa;
    defparam add_223_1.INJECT1_0 = "NO";
    defparam add_223_1.INJECT1_1 = "NO";
    CCU2D add_15371_6 (.A0(addOut[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18717), .COUT(n18718));
    defparam add_15371_6.INIT0 = 16'h5555;
    defparam add_15371_6.INIT1 = 16'h5555;
    defparam add_15371_6.INJECT1_0 = "NO";
    defparam add_15371_6.INJECT1_1 = "NO";
    CCU2D add_15381_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[0]), .B1(speed_set_m1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18609));
    defparam add_15381_1.INIT0 = 16'hF000;
    defparam add_15381_1.INIT1 = 16'ha666;
    defparam add_15381_1.INJECT1_0 = "NO";
    defparam add_15381_1.INJECT1_1 = "NO";
    CCU2D add_15371_4 (.A0(addOut[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18716), .COUT(n18717));
    defparam add_15371_4.INIT0 = 16'h5aaa;
    defparam add_15371_4.INIT1 = 16'h5aaa;
    defparam add_15371_4.INJECT1_0 = "NO";
    defparam add_15371_4.INJECT1_1 = "NO";
    CCU2D add_15371_2 (.A0(addOut[6]), .B0(addOut[5]), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18716));
    defparam add_15371_2.INIT0 = 16'h7000;
    defparam add_15371_2.INIT1 = 16'h5555;
    defparam add_15371_2.INJECT1_0 = "NO";
    defparam add_15371_2.INJECT1_1 = "NO";
    CCU2D add_15372_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18715), 
          .S0(n3780));
    defparam add_15372_cout.INIT0 = 16'h0000;
    defparam add_15372_cout.INIT1 = 16'h0000;
    defparam add_15372_cout.INJECT1_0 = "NO";
    defparam add_15372_cout.INJECT1_1 = "NO";
    CCU2D add_15372_20 (.A0(speed_set_m4[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18714), .COUT(n18715));
    defparam add_15372_20.INIT0 = 16'h5aaa;
    defparam add_15372_20.INIT1 = 16'h0aaa;
    defparam add_15372_20.INJECT1_0 = "NO";
    defparam add_15372_20.INJECT1_1 = "NO";
    CCU2D add_15372_18 (.A0(speed_set_m4[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18713), .COUT(n18714));
    defparam add_15372_18.INIT0 = 16'h5aaa;
    defparam add_15372_18.INIT1 = 16'h5aaa;
    defparam add_15372_18.INJECT1_0 = "NO";
    defparam add_15372_18.INJECT1_1 = "NO";
    CCU2D add_15372_16 (.A0(speed_set_m4[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18712), .COUT(n18713));
    defparam add_15372_16.INIT0 = 16'h5aaa;
    defparam add_15372_16.INIT1 = 16'h5aaa;
    defparam add_15372_16.INJECT1_0 = "NO";
    defparam add_15372_16.INJECT1_1 = "NO";
    CCU2D add_15372_14 (.A0(speed_set_m4[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18711), .COUT(n18712));
    defparam add_15372_14.INIT0 = 16'h5555;
    defparam add_15372_14.INIT1 = 16'h5aaa;
    defparam add_15372_14.INJECT1_0 = "NO";
    defparam add_15372_14.INJECT1_1 = "NO";
    CCU2D add_15372_12 (.A0(speed_set_m4[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18710), .COUT(n18711));
    defparam add_15372_12.INIT0 = 16'h5aaa;
    defparam add_15372_12.INIT1 = 16'h5aaa;
    defparam add_15372_12.INJECT1_0 = "NO";
    defparam add_15372_12.INJECT1_1 = "NO";
    CCU2D add_219_17 (.A0(Out2[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18444), 
          .S0(n1336[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_17.INIT0 = 16'h5aaa;
    defparam add_219_17.INIT1 = 16'h0000;
    defparam add_219_17.INJECT1_0 = "NO";
    defparam add_219_17.INJECT1_1 = "NO";
    CCU2D add_219_15 (.A0(Out2[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18443), 
          .COUT(n18444), .S0(n1336[13]), .S1(n1336[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_15.INIT0 = 16'h5aaa;
    defparam add_219_15.INIT1 = 16'h5aaa;
    defparam add_219_15.INJECT1_0 = "NO";
    defparam add_219_15.INJECT1_1 = "NO";
    CCU2D add_219_13 (.A0(Out2[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18442), 
          .COUT(n18443), .S0(n1336[11]), .S1(n1336[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_13.INIT0 = 16'h5aaa;
    defparam add_219_13.INIT1 = 16'h5aaa;
    defparam add_219_13.INJECT1_0 = "NO";
    defparam add_219_13.INJECT1_1 = "NO";
    CCU2D add_211_9 (.A0(Out0[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18424), 
          .COUT(n18425), .S0(n1294[7]), .S1(n1294[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_9.INIT0 = 16'h5aaa;
    defparam add_211_9.INIT1 = 16'h5aaa;
    defparam add_211_9.INJECT1_0 = "NO";
    defparam add_211_9.INJECT1_1 = "NO";
    CCU2D add_211_7 (.A0(Out0[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18423), 
          .COUT(n18424), .S0(n1294[5]), .S1(n1294[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_7.INIT0 = 16'h5aaa;
    defparam add_211_7.INIT1 = 16'h5aaa;
    defparam add_211_7.INJECT1_0 = "NO";
    defparam add_211_7.INJECT1_1 = "NO";
    CCU2D add_219_11 (.A0(Out2[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18441), 
          .COUT(n18442), .S0(n1336[9]), .S1(n1336[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_11.INIT0 = 16'h5aaa;
    defparam add_219_11.INIT1 = 16'h5aaa;
    defparam add_219_11.INJECT1_0 = "NO";
    defparam add_219_11.INJECT1_1 = "NO";
    CCU2D add_15374_17 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18812), .S1(n3708));
    defparam add_15374_17.INIT0 = 16'h5555;
    defparam add_15374_17.INIT1 = 16'h0000;
    defparam add_15374_17.INJECT1_0 = "NO";
    defparam add_15374_17.INJECT1_1 = "NO";
    CCU2D add_15372_10 (.A0(speed_set_m4[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18709), .COUT(n18710));
    defparam add_15372_10.INIT0 = 16'h5555;
    defparam add_15372_10.INIT1 = 16'h5555;
    defparam add_15372_10.INJECT1_0 = "NO";
    defparam add_15372_10.INJECT1_1 = "NO";
    CCU2D add_15372_8 (.A0(speed_set_m4[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18708), .COUT(n18709));
    defparam add_15372_8.INIT0 = 16'h5aaa;
    defparam add_15372_8.INIT1 = 16'h5555;
    defparam add_15372_8.INJECT1_0 = "NO";
    defparam add_15372_8.INJECT1_1 = "NO";
    CCU2D add_1185_11 (.A0(n1357[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18507), 
          .S0(n2297[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1185_11.INIT0 = 16'hf555;
    defparam add_1185_11.INIT1 = 16'h0000;
    defparam add_1185_11.INJECT1_0 = "NO";
    defparam add_1185_11.INJECT1_1 = "NO";
    CCU2D add_15372_6 (.A0(speed_set_m4[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18707), .COUT(n18708));
    defparam add_15372_6.INIT0 = 16'h5aaa;
    defparam add_15372_6.INIT1 = 16'h5aaa;
    defparam add_15372_6.INJECT1_0 = "NO";
    defparam add_15372_6.INJECT1_1 = "NO";
    CCU2D add_15372_4 (.A0(speed_set_m4[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18706), .COUT(n18707));
    defparam add_15372_4.INIT0 = 16'h5555;
    defparam add_15372_4.INIT1 = 16'h5aaa;
    defparam add_15372_4.INJECT1_0 = "NO";
    defparam add_15372_4.INJECT1_1 = "NO";
    CCU2D add_15374_15 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18811), .COUT(n18812));
    defparam add_15374_15.INIT0 = 16'hf555;
    defparam add_15374_15.INIT1 = 16'hf555;
    defparam add_15374_15.INJECT1_0 = "NO";
    defparam add_15374_15.INJECT1_1 = "NO";
    CCU2D add_15374_13 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18810), .COUT(n18811));
    defparam add_15374_13.INIT0 = 16'hf555;
    defparam add_15374_13.INIT1 = 16'hf555;
    defparam add_15374_13.INJECT1_0 = "NO";
    defparam add_15374_13.INJECT1_1 = "NO";
    CCU2D add_15372_2 (.A0(speed_set_m4[1]), .B0(speed_set_m4[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18706));
    defparam add_15372_2.INIT0 = 16'h1000;
    defparam add_15372_2.INIT1 = 16'h5555;
    defparam add_15372_2.INJECT1_0 = "NO";
    defparam add_15372_2.INJECT1_1 = "NO";
    CCU2D add_1185_9 (.A0(n1357[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1357[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18506), 
          .COUT(n18507), .S0(n2297[7]), .S1(n2297[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1185_9.INIT0 = 16'hf555;
    defparam add_1185_9.INIT1 = 16'hf555;
    defparam add_1185_9.INJECT1_0 = "NO";
    defparam add_1185_9.INJECT1_1 = "NO";
    CCU2D add_15373_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18705), 
          .S0(n3732));
    defparam add_15373_cout.INIT0 = 16'h0000;
    defparam add_15373_cout.INIT1 = 16'h0000;
    defparam add_15373_cout.INJECT1_0 = "NO";
    defparam add_15373_cout.INJECT1_1 = "NO";
    CCU2D add_15373_20 (.A0(speed_set_m3[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18704), .COUT(n18705));
    defparam add_15373_20.INIT0 = 16'h5aaa;
    defparam add_15373_20.INIT1 = 16'h0aaa;
    defparam add_15373_20.INJECT1_0 = "NO";
    defparam add_15373_20.INJECT1_1 = "NO";
    CCU2D add_15373_18 (.A0(speed_set_m3[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18703), .COUT(n18704));
    defparam add_15373_18.INIT0 = 16'h5aaa;
    defparam add_15373_18.INIT1 = 16'h5aaa;
    defparam add_15373_18.INJECT1_0 = "NO";
    defparam add_15373_18.INJECT1_1 = "NO";
    CCU2D add_15374_11 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18809), .COUT(n18810));
    defparam add_15374_11.INIT0 = 16'hf555;
    defparam add_15374_11.INIT1 = 16'hf555;
    defparam add_15374_11.INJECT1_0 = "NO";
    defparam add_15374_11.INJECT1_1 = "NO";
    CCU2D add_15374_9 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18808), .COUT(n18809));
    defparam add_15374_9.INIT0 = 16'hf555;
    defparam add_15374_9.INIT1 = 16'h0aaa;
    defparam add_15374_9.INJECT1_0 = "NO";
    defparam add_15374_9.INJECT1_1 = "NO";
    CCU2D add_15373_16 (.A0(speed_set_m3[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18702), .COUT(n18703));
    defparam add_15373_16.INIT0 = 16'h5aaa;
    defparam add_15373_16.INIT1 = 16'h5aaa;
    defparam add_15373_16.INJECT1_0 = "NO";
    defparam add_15373_16.INJECT1_1 = "NO";
    CCU2D add_15373_14 (.A0(speed_set_m3[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18701), .COUT(n18702));
    defparam add_15373_14.INIT0 = 16'h5555;
    defparam add_15373_14.INIT1 = 16'h5aaa;
    defparam add_15373_14.INJECT1_0 = "NO";
    defparam add_15373_14.INJECT1_1 = "NO";
    CCU2D add_15373_12 (.A0(speed_set_m3[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18700), .COUT(n18701));
    defparam add_15373_12.INIT0 = 16'h5aaa;
    defparam add_15373_12.INIT1 = 16'h5aaa;
    defparam add_15373_12.INJECT1_0 = "NO";
    defparam add_15373_12.INJECT1_1 = "NO";
    CCU2D add_15374_7 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18807), .COUT(n18808));
    defparam add_15374_7.INIT0 = 16'h0aaa;
    defparam add_15374_7.INIT1 = 16'hf555;
    defparam add_15374_7.INJECT1_0 = "NO";
    defparam add_15374_7.INJECT1_1 = "NO";
    CCU2D add_15374_5 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18806), .COUT(n18807));
    defparam add_15374_5.INIT0 = 16'h0aaa;
    defparam add_15374_5.INIT1 = 16'h0aaa;
    defparam add_15374_5.INJECT1_0 = "NO";
    defparam add_15374_5.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_29 (.A0(multOut[27]), .B0(n16283), .C0(addOut[27]), 
          .D0(addIn2_28__N_1440[27]), .A1(multOut[28]), .B1(n16283), .C1(addOut[28]), 
          .D1(addIn2_28__N_1440[28]), .CIN(n18589), .S0(n121[27]), .S1(n121[28]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_29.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_29.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_29.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_29.INJECT1_1 = "NO";
    CCU2D add_1185_7 (.A0(n1357[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1357[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18505), 
          .COUT(n18506), .S0(n2297[5]), .S1(n2297[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1185_7.INIT0 = 16'hf555;
    defparam add_1185_7.INIT1 = 16'hf555;
    defparam add_1185_7.INJECT1_0 = "NO";
    defparam add_1185_7.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_27 (.A0(multOut[25]), .B0(n16283), .C0(addOut[25]), 
          .D0(addIn2_28__N_1440[25]), .A1(multOut[26]), .B1(n16283), .C1(addOut[26]), 
          .D1(addIn2_28__N_1440[26]), .CIN(n18588), .COUT(n18589), .S0(n121[25]), 
          .S1(n121[26]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_27.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_27.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_27.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_27.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_25 (.A0(multOut[23]), .B0(n16283), .C0(addOut[23]), 
          .D0(addIn2_28__N_1440[23]), .A1(multOut[24]), .B1(n16283), .C1(addOut[24]), 
          .D1(addIn2_28__N_1440[24]), .CIN(n18587), .COUT(n18588), .S0(n121[23]), 
          .S1(n121[24]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_25.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_25.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_25.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_25.INJECT1_1 = "NO";
    CCU2D add_15373_10 (.A0(speed_set_m3[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18699), .COUT(n18700));
    defparam add_15373_10.INIT0 = 16'h5555;
    defparam add_15373_10.INIT1 = 16'h5555;
    defparam add_15373_10.INJECT1_0 = "NO";
    defparam add_15373_10.INJECT1_1 = "NO";
    CCU2D add_1185_5 (.A0(n1357[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1357[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18504), 
          .COUT(n18505), .S0(n2297[3]), .S1(n2297[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1185_5.INIT0 = 16'hf555;
    defparam add_1185_5.INIT1 = 16'hf555;
    defparam add_1185_5.INJECT1_0 = "NO";
    defparam add_1185_5.INJECT1_1 = "NO";
    CCU2D add_15374_3 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18805), .COUT(n18806));
    defparam add_15374_3.INIT0 = 16'hf555;
    defparam add_15374_3.INIT1 = 16'hf555;
    defparam add_15374_3.INJECT1_0 = "NO";
    defparam add_15374_3.INJECT1_1 = "NO";
    CCU2D add_15373_8 (.A0(speed_set_m3[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18698), .COUT(n18699));
    defparam add_15373_8.INIT0 = 16'h5aaa;
    defparam add_15373_8.INIT1 = 16'h5555;
    defparam add_15373_8.INJECT1_0 = "NO";
    defparam add_15373_8.INJECT1_1 = "NO";
    FD1P3IX dutyout_m1_i0_i0 (.D(n2261[0]), .SP(clk_N_875_enable_391), .CD(n14336), 
            .CK(clk_N_875), .Q(PWMdut_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i0.GSR = "DISABLED";
    CCU2D addOut_2102_add_4_23 (.A0(multOut[21]), .B0(n16283), .C0(addOut[21]), 
          .D0(addIn2_28__N_1440[21]), .A1(multOut[22]), .B1(n16283), .C1(addOut[22]), 
          .D1(addIn2_28__N_1440[22]), .CIN(n18586), .COUT(n18587), .S0(n121[21]), 
          .S1(n121[22]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_23.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_23.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_23.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_23.INJECT1_1 = "NO";
    CCU2D add_15374_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[4]), .B1(speed_set_m3[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18805));
    defparam add_15374_1.INIT0 = 16'hF000;
    defparam add_15374_1.INIT1 = 16'ha666;
    defparam add_15374_1.INJECT1_0 = "NO";
    defparam add_15374_1.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_21 (.A0(multOut[19]), .B0(n16283), .C0(addOut[19]), 
          .D0(addIn2_28__N_1440[19]), .A1(multOut[20]), .B1(n16283), .C1(addOut[20]), 
          .D1(addIn2_28__N_1440[20]), .CIN(n18585), .COUT(n18586), .S0(n121[19]), 
          .S1(n121[20]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_21.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_21.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_21.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_21.INJECT1_1 = "NO";
    CCU2D add_15373_6 (.A0(speed_set_m3[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18697), .COUT(n18698));
    defparam add_15373_6.INIT0 = 16'h5aaa;
    defparam add_15373_6.INIT1 = 16'h5aaa;
    defparam add_15373_6.INJECT1_0 = "NO";
    defparam add_15373_6.INJECT1_1 = "NO";
    CCU2D add_15375_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18804), 
          .S0(n3684));
    defparam add_15375_cout.INIT0 = 16'h0000;
    defparam add_15375_cout.INIT1 = 16'h0000;
    defparam add_15375_cout.INJECT1_0 = "NO";
    defparam add_15375_cout.INJECT1_1 = "NO";
    CCU2D add_219_9 (.A0(Out2[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18440), 
          .COUT(n18441), .S0(n1336[7]), .S1(n1336[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_9.INIT0 = 16'h5aaa;
    defparam add_219_9.INIT1 = 16'h5aaa;
    defparam add_219_9.INJECT1_0 = "NO";
    defparam add_219_9.INJECT1_1 = "NO";
    LUT4 mux_1253_i8_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[7]), 
         .D(speed_set_m4[7]), .Z(n2593[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i8_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1185_3 (.A0(n1357[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1357[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18503), 
          .COUT(n18504), .S0(n2297[1]), .S1(n2297[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1185_3.INIT0 = 16'hf555;
    defparam add_1185_3.INIT1 = 16'hf555;
    defparam add_1185_3.INJECT1_0 = "NO";
    defparam add_1185_3.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_19 (.A0(multOut[17]), .B0(n16283), .C0(addOut[17]), 
          .D0(addIn2_28__N_1440[17]), .A1(multOut[18]), .B1(n16283), .C1(addOut[18]), 
          .D1(addIn2_28__N_1440[18]), .CIN(n18584), .COUT(n18585), .S0(n121[17]), 
          .S1(n121[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_19.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_19.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_19.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_19.INJECT1_1 = "NO";
    CCU2D add_219_7 (.A0(Out2[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18439), 
          .COUT(n18440), .S0(n1336[5]), .S1(n1336[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_7.INIT0 = 16'h5aaa;
    defparam add_219_7.INIT1 = 16'h5aaa;
    defparam add_219_7.INJECT1_0 = "NO";
    defparam add_219_7.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_17 (.A0(multOut[15]), .B0(n16283), .C0(addOut[15]), 
          .D0(addIn2_28__N_1440[15]), .A1(multOut[16]), .B1(n16283), .C1(addOut[16]), 
          .D1(addIn2_28__N_1440[16]), .CIN(n18583), .COUT(n18584), .S0(n121[15]), 
          .S1(n121[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_17.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_17.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_17.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_17.INJECT1_1 = "NO";
    CCU2D add_15373_4 (.A0(speed_set_m3[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18696), .COUT(n18697));
    defparam add_15373_4.INIT0 = 16'h5555;
    defparam add_15373_4.INIT1 = 16'h5aaa;
    defparam add_15373_4.INJECT1_0 = "NO";
    defparam add_15373_4.INJECT1_1 = "NO";
    CCU2D add_219_5 (.A0(Out2[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18438), 
          .COUT(n18439), .S0(n1336[3]), .S1(n1336[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_5.INIT0 = 16'h5aaa;
    defparam add_219_5.INIT1 = 16'h5aaa;
    defparam add_219_5.INJECT1_0 = "NO";
    defparam add_219_5.INJECT1_1 = "NO";
    CCU2D add_1185_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1357[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18503), 
          .S1(n2297[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1185_1.INIT0 = 16'hF000;
    defparam add_1185_1.INIT1 = 16'h0aaa;
    defparam add_1185_1.INJECT1_0 = "NO";
    defparam add_1185_1.INJECT1_1 = "NO";
    CCU2D add_15373_2 (.A0(speed_set_m3[1]), .B0(speed_set_m3[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18696));
    defparam add_15373_2.INIT0 = 16'h1000;
    defparam add_15373_2.INIT1 = 16'h5555;
    defparam add_15373_2.INJECT1_0 = "NO";
    defparam add_15373_2.INJECT1_1 = "NO";
    CCU2D add_15375_20 (.A0(speed_set_m2[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18803), .COUT(n18804));
    defparam add_15375_20.INIT0 = 16'h5aaa;
    defparam add_15375_20.INIT1 = 16'h0aaa;
    defparam add_15375_20.INJECT1_0 = "NO";
    defparam add_15375_20.INJECT1_1 = "NO";
    CCU2D add_15375_18 (.A0(speed_set_m2[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18802), .COUT(n18803));
    defparam add_15375_18.INIT0 = 16'h5aaa;
    defparam add_15375_18.INIT1 = 16'h5aaa;
    defparam add_15375_18.INJECT1_0 = "NO";
    defparam add_15375_18.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_15 (.A0(multOut[13]), .B0(n16283), .C0(addOut[13]), 
          .D0(addIn2_28__N_1440[13]), .A1(multOut[14]), .B1(n16283), .C1(addOut[14]), 
          .D1(addIn2_28__N_1440[14]), .CIN(n18582), .COUT(n18583), .S0(n121[13]), 
          .S1(n121[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_15.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_15.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_15.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_15.INJECT1_1 = "NO";
    LUT4 i1755_1_lut (.A(n42), .Z(subIn1_24__N_1533)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(137[34:50])
    defparam i1755_1_lut.init = 16'h5555;
    CCU2D add_211_5 (.A0(Out0[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18422), 
          .COUT(n18423), .S0(n1294[3]), .S1(n1294[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_5.INIT0 = 16'h5aaa;
    defparam add_211_5.INIT1 = 16'h5aaa;
    defparam add_211_5.INJECT1_0 = "NO";
    defparam add_211_5.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_13 (.A0(multOut[11]), .B0(n16283), .C0(addOut[11]), 
          .D0(addIn2_28__N_1440[11]), .A1(multOut[12]), .B1(n16283), .C1(addOut[12]), 
          .D1(addIn2_28__N_1440[12]), .CIN(n18581), .COUT(n18582), .S0(n121[11]), 
          .S1(n121[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_13.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_13.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_13.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_13.INJECT1_1 = "NO";
    CCU2D add_15375_16 (.A0(speed_set_m2[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18801), .COUT(n18802));
    defparam add_15375_16.INIT0 = 16'h5aaa;
    defparam add_15375_16.INIT1 = 16'h5aaa;
    defparam add_15375_16.INJECT1_0 = "NO";
    defparam add_15375_16.INJECT1_1 = "NO";
    LUT4 i1756_1_lut (.A(n49), .Z(dirout_m3_N_1947)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(139[35:51])
    defparam i1756_1_lut.init = 16'h5555;
    LUT4 i1754_1_lut (.A(n35), .Z(subIn1_24__N_1347)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(135[34:50])
    defparam i1754_1_lut.init = 16'h5555;
    CCU2D addOut_2102_add_4_11 (.A0(multOut[9]), .B0(n16283), .C0(addOut[9]), 
          .D0(addIn2_28__N_1440[9]), .A1(multOut[10]), .B1(n16283), .C1(addOut[10]), 
          .D1(addIn2_28__N_1440[10]), .CIN(n18580), .COUT(n18581), .S0(n121[9]), 
          .S1(n121[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_11.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_11.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_11.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_11.INJECT1_1 = "NO";
    CCU2D add_15375_14 (.A0(speed_set_m2[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18800), .COUT(n18801));
    defparam add_15375_14.INIT0 = 16'h5555;
    defparam add_15375_14.INIT1 = 16'h5aaa;
    defparam add_15375_14.INJECT1_0 = "NO";
    defparam add_15375_14.INJECT1_1 = "NO";
    LUT4 mux_1253_i12_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[11]), 
         .D(speed_set_m4[11]), .Z(n2593[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i12_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15375_12 (.A0(speed_set_m2[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18799), .COUT(n18800));
    defparam add_15375_12.INIT0 = 16'h5aaa;
    defparam add_15375_12.INIT1 = 16'h5aaa;
    defparam add_15375_12.INJECT1_0 = "NO";
    defparam add_15375_12.INJECT1_1 = "NO";
    LUT4 i1757_1_lut (.A(n56), .Z(dirout_m4_N_1950)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(141[35:51])
    defparam i1757_1_lut.init = 16'h5555;
    CCU2D add_1184_11 (.A0(n1336[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18502), 
          .S0(n2285[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1184_11.INIT0 = 16'hf555;
    defparam add_1184_11.INIT1 = 16'h0000;
    defparam add_1184_11.INJECT1_0 = "NO";
    defparam add_1184_11.INJECT1_1 = "NO";
    CCU2D add_1184_9 (.A0(n1336[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1336[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18501), 
          .COUT(n18502), .S0(n2285[7]), .S1(n2285[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1184_9.INIT0 = 16'hf555;
    defparam add_1184_9.INIT1 = 16'hf555;
    defparam add_1184_9.INJECT1_0 = "NO";
    defparam add_1184_9.INJECT1_1 = "NO";
    LUT4 mux_1253_i13_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[12]), 
         .D(speed_set_m4[12]), .Z(n2593[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13364_2_lut (.A(addOut[28]), .B(n22440), .Z(Out0_28__N_1087[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13364_2_lut.init = 16'h2222;
    CCU2D addOut_2102_add_4_9 (.A0(multOut[7]), .B0(n16283), .C0(addOut[7]), 
          .D0(addIn2_28__N_1440[7]), .A1(multOut[8]), .B1(n16283), .C1(addOut[8]), 
          .D1(addIn2_28__N_1440[8]), .CIN(n18579), .COUT(n18580), .S0(n121[7]), 
          .S1(n121[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_9.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_9.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_9.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_9.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_7 (.A0(multOut[5]), .B0(n16283), .C0(addOut[5]), 
          .D0(addIn2_28__N_1440[5]), .A1(multOut[6]), .B1(n16283), .C1(addOut[6]), 
          .D1(addIn2_28__N_1440[6]), .CIN(n18578), .COUT(n18579), .S0(n121[5]), 
          .S1(n121[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_7.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_7.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_7.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_7.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_5 (.A0(multOut[3]), .B0(n16283), .C0(addOut[3]), 
          .D0(addIn2_28__N_1440[3]), .A1(multOut[4]), .B1(n16283), .C1(addOut[4]), 
          .D1(addIn2_28__N_1440[4]), .CIN(n18577), .COUT(n18578), .S0(n121[3]), 
          .S1(n121[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_5.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_5.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_5.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_5.INJECT1_1 = "NO";
    LUT4 mux_1253_i14_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[13]), 
         .D(speed_set_m4[13]), .Z(n2593[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i14_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15375_10 (.A0(speed_set_m2[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18798), .COUT(n18799));
    defparam add_15375_10.INIT0 = 16'h5555;
    defparam add_15375_10.INIT1 = 16'h5555;
    defparam add_15375_10.INJECT1_0 = "NO";
    defparam add_15375_10.INJECT1_1 = "NO";
    CCU2D add_15375_8 (.A0(speed_set_m2[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18797), .COUT(n18798));
    defparam add_15375_8.INIT0 = 16'h5aaa;
    defparam add_15375_8.INIT1 = 16'h5555;
    defparam add_15375_8.INJECT1_0 = "NO";
    defparam add_15375_8.INJECT1_1 = "NO";
    CCU2D add_1184_7 (.A0(n1336[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1336[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18500), 
          .COUT(n18501), .S0(n2285[5]), .S1(n2285[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1184_7.INIT0 = 16'hf555;
    defparam add_1184_7.INIT1 = 16'hf555;
    defparam add_1184_7.INJECT1_0 = "NO";
    defparam add_1184_7.INJECT1_1 = "NO";
    LUT4 i13359_2_lut (.A(addOut[27]), .B(n22440), .Z(Out0_28__N_1087[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13359_2_lut.init = 16'h2222;
    LUT4 i7_4_lut_adj_105 (.A(Out2[3]), .B(n14_adj_2366), .C(n10_adj_2367), 
         .D(Out2[4]), .Z(n18892)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i7_4_lut_adj_105.init = 16'hfffe;
    CCU2D add_1184_5 (.A0(n1336[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1336[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18499), 
          .COUT(n18500), .S0(n2285[3]), .S1(n2285[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1184_5.INIT0 = 16'hf555;
    defparam add_1184_5.INIT1 = 16'hf555;
    defparam add_1184_5.INJECT1_0 = "NO";
    defparam add_1184_5.INJECT1_1 = "NO";
    CCU2D addOut_2102_add_4_3 (.A0(multOut[1]), .B0(n16283), .C0(addOut[1]), 
          .D0(addIn2_28__N_1440[1]), .A1(multOut[2]), .B1(n16283), .C1(addOut[2]), 
          .D1(addIn2_28__N_1440[2]), .CIN(n18576), .COUT(n18577), .S0(n121[1]), 
          .S1(n121[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_3.INIT0 = 16'h569a;
    defparam addOut_2102_add_4_3.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_3.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_3.INJECT1_1 = "NO";
    LUT4 i6_4_lut_adj_106 (.A(Out2[11]), .B(Out2[7]), .C(Out2[2]), .D(Out2[10]), 
         .Z(n14_adj_2366)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i6_4_lut_adj_106.init = 16'hfffe;
    CCU2D addOut_2102_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(multOut[0]), .B1(n16283), .C1(addOut[0]), 
          .D1(addIn2_28__N_1440[0]), .COUT(n18576), .S1(n121[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102_add_4_1.INIT0 = 16'hF000;
    defparam addOut_2102_add_4_1.INIT1 = 16'h569a;
    defparam addOut_2102_add_4_1.INJECT1_0 = "NO";
    defparam addOut_2102_add_4_1.INJECT1_1 = "NO";
    LUT4 i2_2_lut_adj_107 (.A(Out2[9]), .B(Out2[1]), .Z(n10_adj_2367)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i2_2_lut_adj_107.init = 16'heeee;
    CCU2D add_15376_17 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18687), .S1(n3660));
    defparam add_15376_17.INIT0 = 16'h5555;
    defparam add_15376_17.INIT1 = 16'h0000;
    defparam add_15376_17.INJECT1_0 = "NO";
    defparam add_15376_17.INJECT1_1 = "NO";
    PFUMX mux_1202_i21 (.BLUT(n5402), .ALUT(n5360), .C0(n2545), .Z(n5450));
    CCU2D add_15376_15 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18686), .COUT(n18687));
    defparam add_15376_15.INIT0 = 16'hf555;
    defparam add_15376_15.INIT1 = 16'hf555;
    defparam add_15376_15.INJECT1_0 = "NO";
    defparam add_15376_15.INJECT1_1 = "NO";
    PFUMX mux_1202_i20 (.BLUT(n5400), .ALUT(n5358), .C0(n2545), .Z(n5448));
    PFUMX mux_1202_i19 (.BLUT(n5398), .ALUT(n5356), .C0(n2545), .Z(n5446));
    PFUMX mux_1202_i18 (.BLUT(n5396), .ALUT(n5354), .C0(n2545), .Z(n5444));
    PFUMX mux_1202_i17 (.BLUT(n5394), .ALUT(n5352), .C0(n2545), .Z(n5442));
    LUT4 i4_4_lut_adj_108 (.A(Out2[5]), .B(Out2[6]), .C(Out2[0]), .D(n6_adj_2368), 
         .Z(n18893)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i4_4_lut_adj_108.init = 16'hfffe;
    CCU2D add_15376_13 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18685), .COUT(n18686));
    defparam add_15376_13.INIT0 = 16'hf555;
    defparam add_15376_13.INIT1 = 16'hf555;
    defparam add_15376_13.INJECT1_0 = "NO";
    defparam add_15376_13.INJECT1_1 = "NO";
    PFUMX mux_1202_i16 (.BLUT(n5392), .ALUT(n5350), .C0(n2545), .Z(n5440));
    PFUMX mux_1202_i15 (.BLUT(n5390), .ALUT(n5348), .C0(n2545), .Z(n5438));
    PFUMX mux_1202_i14 (.BLUT(n5388), .ALUT(n5346), .C0(n2545), .Z(n5436));
    CCU2D add_15376_11 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18684), .COUT(n18685));
    defparam add_15376_11.INIT0 = 16'hf555;
    defparam add_15376_11.INIT1 = 16'hf555;
    defparam add_15376_11.INJECT1_0 = "NO";
    defparam add_15376_11.INJECT1_1 = "NO";
    PFUMX mux_1202_i13 (.BLUT(n5386), .ALUT(n5344), .C0(n2545), .Z(n5434));
    PFUMX mux_1202_i12 (.BLUT(n5384), .ALUT(n5342), .C0(n2545), .Z(n5432));
    PFUMX mux_1202_i11 (.BLUT(n5382), .ALUT(n5340), .C0(n2545), .Z(n5430));
    PFUMX mux_1202_i10 (.BLUT(n5380), .ALUT(n5338), .C0(n2545), .Z(n5428));
    PFUMX mux_1202_i9 (.BLUT(n5378), .ALUT(n5336), .C0(n2545), .Z(n5426));
    CCU2D add_15375_6 (.A0(speed_set_m2[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18796), .COUT(n18797));
    defparam add_15375_6.INIT0 = 16'h5aaa;
    defparam add_15375_6.INIT1 = 16'h5aaa;
    defparam add_15375_6.INJECT1_0 = "NO";
    defparam add_15375_6.INJECT1_1 = "NO";
    PFUMX mux_1202_i8 (.BLUT(n5376), .ALUT(n5334), .C0(n2545), .Z(n5424));
    PFUMX mux_1202_i7 (.BLUT(n5374), .ALUT(n5332), .C0(n2545), .Z(n5422));
    PFUMX mux_1202_i6 (.BLUT(n5372), .ALUT(n5330), .C0(n2545), .Z(n5420));
    PFUMX mux_1202_i5 (.BLUT(n5370), .ALUT(n5328), .C0(n2545), .Z(n5418));
    CCU2D add_15375_4 (.A0(speed_set_m2[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18795), .COUT(n18796));
    defparam add_15375_4.INIT0 = 16'h5555;
    defparam add_15375_4.INIT1 = 16'h5aaa;
    defparam add_15375_4.INJECT1_0 = "NO";
    defparam add_15375_4.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_109 (.A(Out2[8]), .B(Out2[12]), .Z(n6_adj_2368)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i1_2_lut_adj_109.init = 16'heeee;
    LUT4 i2967_2_lut_rep_380 (.A(n22440), .B(n22435), .Z(clk_N_875_enable_391)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i2967_2_lut_rep_380.init = 16'h8888;
    PFUMX mux_1202_i4 (.BLUT(n5368), .ALUT(n5326), .C0(n2545), .Z(n5416));
    LUT4 i11783_2_lut_3_lut_4_lut (.A(n22440), .B(n22435), .C(n21697), 
         .D(n21698), .Z(n14340)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11783_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 mux_1253_i17_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[16]), 
         .D(speed_set_m4[16]), .Z(n2593[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i17_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_rep_381 (.A(ss[1]), .B(ss[2]), .Z(n21694)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_381.init = 16'h8888;
    PFUMX mux_1202_i3 (.BLUT(n5366), .ALUT(n5324), .C0(n2545), .Z(n5414));
    LUT4 i1_2_lut_rep_363_3_lut (.A(ss[1]), .B(ss[2]), .C(ss[0]), .Z(n21676)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_363_3_lut.init = 16'h8080;
    LUT4 i13284_2_lut (.A(addOut[26]), .B(n22440), .Z(backOut3_28__N_1872[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13284_2_lut.init = 16'h2222;
    CCU2D add_15375_2 (.A0(speed_set_m2[1]), .B0(speed_set_m2[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18795));
    defparam add_15375_2.INIT0 = 16'h1000;
    defparam add_15375_2.INIT1 = 16'h5555;
    defparam add_15375_2.INJECT1_0 = "NO";
    defparam add_15375_2.INJECT1_1 = "NO";
    LUT4 i9146_2_lut_3_lut_4_lut (.A(ss[1]), .B(ss[2]), .C(ss[3]), .D(ss[0]), 
         .Z(n15)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i9146_2_lut_3_lut_4_lut.init = 16'h78f0;
    PFUMX mux_1202_i2 (.BLUT(n5364), .ALUT(n5322), .C0(n2545), .Z(n5412));
    PFUMX mux_1202_i1 (.BLUT(n5320), .ALUT(n5318), .C0(n2545), .Z(n5410));
    LUT4 i1_2_lut_rep_384 (.A(n22433), .B(ss[1]), .Z(n21697)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_384.init = 16'heeee;
    LUT4 i13345_2_lut (.A(addOut[25]), .B(n22440), .Z(Out0_28__N_1087[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13345_2_lut.init = 16'h2222;
    LUT4 i13280_2_lut (.A(addOut[24]), .B(n22440), .Z(backOut3_28__N_1872[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13280_2_lut.init = 16'h2222;
    PFUMX i3024 (.BLUT(n2593[0]), .ALUT(n5518), .C0(n21630), .Z(n5519));
    PFUMX i3311 (.BLUT(n2593[1]), .ALUT(n5805), .C0(n21630), .Z(n5806));
    PFUMX i3313 (.BLUT(n2593[2]), .ALUT(n5807), .C0(n21630), .Z(n5808));
    PFUMX i3315 (.BLUT(n2593[3]), .ALUT(n5809), .C0(n21630), .Z(n5810));
    LUT4 i1_3_lut_rep_361_4_lut (.A(ss[2]), .B(ss[1]), .C(ss[3]), .D(n22440), 
         .Z(n21674)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i1_3_lut_rep_361_4_lut.init = 16'h001e;
    LUT4 i13103_3_lut_4_lut (.A(n21659), .B(n21648), .C(n21658), .D(n21660), 
         .Z(multIn2[8])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;
    defparam i13103_3_lut_4_lut.init = 16'h00f7;
    PFUMX i3317 (.BLUT(n2593[4]), .ALUT(n5811), .C0(n21630), .Z(n5812));
    LUT4 i2_3_lut_4_lut_adj_110 (.A(n22433), .B(ss[1]), .C(ss[3]), .D(ss[0]), 
         .Z(n18943)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_110.init = 16'hfffe;
    PFUMX i3319 (.BLUT(n2593[5]), .ALUT(n5813), .C0(n21630), .Z(n5814));
    PFUMX i3321 (.BLUT(n2593[6]), .ALUT(n5815), .C0(n21630), .Z(n5816));
    LUT4 i1_2_lut_rep_385 (.A(ss[0]), .B(ss[3]), .Z(n21698)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_385.init = 16'heeee;
    LUT4 i3_2_lut_rep_364_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), 
         .D(n22433), .Z(n21677)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i3_2_lut_rep_364_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_91_i13_3_lut_4_lut_4_lut (.A(n21646), .B(\speed_avg_m4[12] ), 
         .C(n4358), .D(n21648), .Z(n367[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i13_3_lut_4_lut_4_lut.init = 16'hcacf;
    PFUMX i3323 (.BLUT(n2593[7]), .ALUT(n5817), .C0(n21630), .Z(n5818));
    CCU2D add_15376_9 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18683), .COUT(n18684));
    defparam add_15376_9.INIT0 = 16'hf555;
    defparam add_15376_9.INIT1 = 16'h0aaa;
    defparam add_15376_9.INJECT1_0 = "NO";
    defparam add_15376_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_111 (.A(ss[0]), .B(ss[3]), .C(n22433), 
         .D(ss[1]), .Z(n19913)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut_4_lut_adj_111.init = 16'h1000;
    CCU2D add_15376_7 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18682), .COUT(n18683));
    defparam add_15376_7.INIT0 = 16'h0aaa;
    defparam add_15376_7.INIT1 = 16'hf555;
    defparam add_15376_7.INJECT1_0 = "NO";
    defparam add_15376_7.INJECT1_1 = "NO";
    PFUMX i3325 (.BLUT(n2593[8]), .ALUT(n5819), .C0(n21630), .Z(n5820));
    LUT4 mux_91_i10_3_lut_4_lut_4_lut (.A(n21646), .B(\speed_avg_m4[9] ), 
         .C(n4358), .D(n21648), .Z(n367[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i10_3_lut_4_lut_4_lut.init = 16'hcacf;
    CCU2D add_1184_3 (.A0(n1336[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1336[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18498), 
          .COUT(n18499), .S0(n2285[1]), .S1(n2285[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1184_3.INIT0 = 16'hf555;
    defparam add_1184_3.INIT1 = 16'hf555;
    defparam add_1184_3.INJECT1_0 = "NO";
    defparam add_1184_3.INJECT1_1 = "NO";
    CCU2D add_1184_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1336[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18498), 
          .S1(n2285[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1184_1.INIT0 = 16'hF000;
    defparam add_1184_1.INIT1 = 16'h0aaa;
    defparam add_1184_1.INJECT1_0 = "NO";
    defparam add_1184_1.INJECT1_1 = "NO";
    CCU2D add_15376_5 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18681), .COUT(n18682));
    defparam add_15376_5.INIT0 = 16'h0aaa;
    defparam add_15376_5.INIT1 = 16'h0aaa;
    defparam add_15376_5.INJECT1_0 = "NO";
    defparam add_15376_5.INJECT1_1 = "NO";
    PFUMX i3327 (.BLUT(n2593[9]), .ALUT(n5821), .C0(n21630), .Z(n5822));
    CCU2D add_15376_3 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18680), .COUT(n18681));
    defparam add_15376_3.INIT0 = 16'hf555;
    defparam add_15376_3.INIT1 = 16'hf555;
    defparam add_15376_3.INJECT1_0 = "NO";
    defparam add_15376_3.INJECT1_1 = "NO";
    LUT4 i2_2_lut_rep_365_3_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n21678)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_2_lut_rep_365_3_lut.init = 16'hefef;
    LUT4 i13566_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), .D(n22433), 
         .Z(n16131)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13566_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 mux_1253_i18_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[17]), 
         .D(speed_set_m4[17]), .Z(n2593[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i18_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_91_i9_3_lut_4_lut_4_lut (.A(n21646), .B(\speed_avg_m4[8] ), 
         .C(n4358), .D(n21648), .Z(n367[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i9_3_lut_4_lut_4_lut.init = 16'hcacf;
    PFUMX i3329 (.BLUT(n2593[10]), .ALUT(n5823), .C0(n21630), .Z(n5824));
    CCU2D add_211_3 (.A0(Out0[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18421), 
          .COUT(n18422), .S0(n1294[1]), .S1(n1294[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_3.INIT0 = 16'h5aaa;
    defparam add_211_3.INIT1 = 16'h5aaa;
    defparam add_211_3.INJECT1_0 = "NO";
    defparam add_211_3.INJECT1_1 = "NO";
    LUT4 mux_91_i8_3_lut_4_lut_4_lut (.A(n21646), .B(\speed_avg_m4[7] ), 
         .C(n4358), .D(n21648), .Z(n367[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i8_3_lut_4_lut_4_lut.init = 16'hcacf;
    PFUMX i3331 (.BLUT(n2593[11]), .ALUT(n5825), .C0(n21630), .Z(n5826));
    LUT4 mux_91_i4_3_lut_4_lut_4_lut (.A(n21646), .B(\speed_avg_m4[3] ), 
         .C(n4358), .D(n21648), .Z(n367[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i4_3_lut_4_lut_4_lut.init = 16'hcacf;
    PFUMX i3333 (.BLUT(n2593[12]), .ALUT(n5827), .C0(n21630), .Z(n5828));
    PFUMX i3335 (.BLUT(n2593[13]), .ALUT(n5829), .C0(n21630), .Z(n5830));
    PFUMX i3337 (.BLUT(n2593[14]), .ALUT(n5831), .C0(n21630), .Z(n5832));
    PFUMX i3339 (.BLUT(n2593[15]), .ALUT(n5833), .C0(n21630), .Z(n5834));
    CCU2D add_1183_11 (.A0(n1315[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18497), 
          .S0(n2273[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1183_11.INIT0 = 16'hf555;
    defparam add_1183_11.INIT1 = 16'h0000;
    defparam add_1183_11.INJECT1_0 = "NO";
    defparam add_1183_11.INJECT1_1 = "NO";
    LUT4 mux_1253_i19_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[18]), 
         .D(speed_set_m4[18]), .Z(n2593[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i19_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1183_9 (.A0(n1315[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1315[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18496), 
          .COUT(n18497), .S0(n2273[7]), .S1(n2273[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1183_9.INIT0 = 16'hf555;
    defparam add_1183_9.INIT1 = 16'hf555;
    defparam add_1183_9.INJECT1_0 = "NO";
    defparam add_1183_9.INJECT1_1 = "NO";
    CCU2D add_15376_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[4]), .B1(speed_set_m2[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18680));
    defparam add_15376_1.INIT0 = 16'hF000;
    defparam add_15376_1.INIT1 = 16'ha666;
    defparam add_15376_1.INJECT1_0 = "NO";
    defparam add_15376_1.INJECT1_1 = "NO";
    LUT4 mux_1253_i20_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[19]), 
         .D(speed_set_m4[19]), .Z(n2593[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i20_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1183_7 (.A0(n1315[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1315[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18495), 
          .COUT(n18496), .S0(n2273[5]), .S1(n2273[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1183_7.INIT0 = 16'hf555;
    defparam add_1183_7.INIT1 = 16'hf555;
    defparam add_1183_7.INJECT1_0 = "NO";
    defparam add_1183_7.INJECT1_1 = "NO";
    CCU2D add_1183_5 (.A0(n1315[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1315[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18494), 
          .COUT(n18495), .S0(n2273[3]), .S1(n2273[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1183_5.INIT0 = 16'hf555;
    defparam add_1183_5.INIT1 = 16'hf555;
    defparam add_1183_5.INJECT1_0 = "NO";
    defparam add_1183_5.INJECT1_1 = "NO";
    CCU2D add_219_3 (.A0(Out2[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18437), 
          .COUT(n18438), .S0(n1336[1]), .S1(n1336[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_3.INIT0 = 16'h5aaa;
    defparam add_219_3.INIT1 = 16'h5aaa;
    defparam add_219_3.INJECT1_0 = "NO";
    defparam add_219_3.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_23 (.A0(n8_adj_2369), .B0(n16337), .C0(n5846), 
          .D0(n16073), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18679), .S0(n4479));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_23.INIT0 = 16'h0f8f;
    defparam sub_16_rep_4_add_2_23.INIT1 = 16'h0000;
    defparam sub_16_rep_4_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_23.INJECT1_1 = "NO";
    PFUMX i3341 (.BLUT(n2593[16]), .ALUT(n5835), .C0(n21630), .Z(n5836));
    PFUMX i3343 (.BLUT(n2593[17]), .ALUT(n5837), .C0(n21630), .Z(n5838));
    CCU2D add_219_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[13]), .B1(n18892), .C1(n18893), .D1(Out2[28]), .COUT(n18437), 
          .S1(n1336[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_1.INIT0 = 16'hF000;
    defparam add_219_1.INIT1 = 16'h56aa;
    defparam add_219_1.INJECT1_0 = "NO";
    defparam add_219_1.INJECT1_1 = "NO";
    PFUMX i3345 (.BLUT(n2593[18]), .ALUT(n5839), .C0(n21630), .Z(n5840));
    PFUMX i3347 (.BLUT(n2593[19]), .ALUT(n5841), .C0(n21630), .Z(n5842));
    PFUMX i3351 (.BLUT(n2593[20]), .ALUT(n5845), .C0(n21630), .Z(n5846));
    L6MUX21 addIn2_28__I_29_i25 (.D0(n615[24]), .D1(addIn2_28__N_1569[24]), 
            .SD(n20384), .Z(addIn2_28__N_1440[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13341_2_lut (.A(addOut[23]), .B(n22440), .Z(Out0_28__N_1087[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13341_2_lut.init = 16'h2222;
    L6MUX21 addIn2_28__I_29_i4 (.D0(n615[3]), .D1(addIn2_28__N_1569[3]), 
            .SD(n20384), .Z(addIn2_28__N_1440[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_1183_3 (.A0(n1315[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1315[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18493), 
          .COUT(n18494), .S0(n2273[1]), .S1(n2273[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1183_3.INIT0 = 16'hf555;
    defparam add_1183_3.INIT1 = 16'hf555;
    defparam add_1183_3.INJECT1_0 = "NO";
    defparam add_1183_3.INJECT1_1 = "NO";
    L6MUX21 addIn2_28__I_29_i26 (.D0(n615[25]), .D1(addIn2_28__N_1569[25]), 
            .SD(n20384), .Z(addIn2_28__N_1440[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i5 (.D0(n615[4]), .D1(addIn2_28__N_1569[4]), 
            .SD(n20384), .Z(addIn2_28__N_1440[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i27 (.D0(n615[26]), .D1(addIn2_28__N_1569[26]), 
            .SD(n20384), .Z(addIn2_28__N_1440[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i6 (.D0(n615[5]), .D1(addIn2_28__N_1569[5]), 
            .SD(n20384), .Z(addIn2_28__N_1440[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D sub_16_rep_4_add_2_21 (.A0(n4409), .B0(n11474), .C0(n5842), 
          .D0(n16073), .A1(n8_adj_2369), .B1(n16337), .C1(n5846), .D1(n16073), 
          .CIN(n18678), .COUT(n18679), .S0(n4481), .S1(n4480));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_21.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_21.INIT1 = 16'h0f8f;
    defparam sub_16_rep_4_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_19 (.A0(n4411), .B0(n11474), .C0(n5838), 
          .D0(n16073), .A1(n4410), .B1(n11474), .C1(n5840), .D1(n16073), 
          .CIN(n18677), .COUT(n18678), .S0(n4483), .S1(n4482));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_19.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_19.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_19.INJECT1_1 = "NO";
    FD1P3IX dutyout_m4_i0_i9 (.D(n19337), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i8 (.D(n19331), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i7 (.D(n19325), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i6 (.D(n1539[6]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i6.GSR = "DISABLED";
    CCU2D sub_16_rep_4_add_2_17 (.A0(n4413), .B0(n11474), .C0(n5834), 
          .D0(n16073), .A1(n4412), .B1(n11474), .C1(n5836), .D1(n16073), 
          .CIN(n18676), .COUT(n18677), .S0(n4485), .S1(n4484));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_17.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_17.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_17.INJECT1_1 = "NO";
    CCU2D add_1183_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1315[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18493), 
          .S1(n2273[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1183_1.INIT0 = 16'hF000;
    defparam add_1183_1.INIT1 = 16'h0aaa;
    defparam add_1183_1.INJECT1_0 = "NO";
    defparam add_1183_1.INJECT1_1 = "NO";
    FD1P3IX dutyout_m4_i0_i5 (.D(n1539[5]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i4 (.D(n2297[4]), .SP(clk_N_875_enable_391), .CD(n14363), 
            .CK(clk_N_875), .Q(PWMdut_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i3 (.D(n1539[3]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i2 (.D(n2297[2]), .SP(clk_N_875_enable_391), .CD(n14363), 
            .CK(clk_N_875), .Q(PWMdut_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i1 (.D(n2297[1]), .SP(clk_N_875_enable_391), .CD(n14363), 
            .CK(clk_N_875), .Q(PWMdut_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i9 (.D(n1495[9]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i8 (.D(n1495[8]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i8.GSR = "DISABLED";
    CCU2D sub_16_rep_4_add_2_15 (.A0(n4415), .B0(n11474), .C0(n5830), 
          .D0(n16073), .A1(n4414), .B1(n11474), .C1(n5832), .D1(n16073), 
          .CIN(n18675), .COUT(n18676), .S0(n4487), .S1(n4486));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_15.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_15.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_15.INJECT1_1 = "NO";
    FD1P3IX dutyout_m3_i0_i7 (.D(n1495[7]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i6 (.D(n1495[6]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i5 (.D(n1495[5]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i4 (.D(n2285[4]), .SP(clk_N_875_enable_391), .CD(n14354), 
            .CK(clk_N_875), .Q(PWMdut_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i3 (.D(n1495[3]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i2 (.D(n2285[2]), .SP(clk_N_875_enable_391), .CD(n14354), 
            .CK(clk_N_875), .Q(PWMdut_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i1 (.D(n2285[1]), .SP(clk_N_875_enable_391), .CD(n14354), 
            .CK(clk_N_875), .Q(PWMdut_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i9 (.D(n19319), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i8 (.D(n19313), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i7 (.D(n19307), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i6 (.D(n1451[6]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i5 (.D(n1451[5]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i4 (.D(n2273[4]), .SP(clk_N_875_enable_391), .CD(n14345), 
            .CK(clk_N_875), .Q(PWMdut_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i3 (.D(n1451[3]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i2 (.D(n2273[2]), .SP(clk_N_875_enable_391), .CD(n14345), 
            .CK(clk_N_875), .Q(PWMdut_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i1 (.D(n2273[1]), .SP(clk_N_875_enable_391), .CD(n14345), 
            .CK(clk_N_875), .Q(PWMdut_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i9 (.D(n1407[9]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i8 (.D(n1407[8]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i7 (.D(n1407[7]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i6 (.D(n1407[6]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i6.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i28 (.D0(n615[27]), .D1(addIn2_28__N_1569[27]), 
            .SD(n20384), .Z(addIn2_28__N_1440[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX dutyout_m1_i0_i5 (.D(n1407[5]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i4 (.D(n2261[4]), .SP(clk_N_875_enable_391), .CD(n14336), 
            .CK(clk_N_875), .Q(PWMdut_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i3 (.D(n1407[3]), .SP(clk_N_875_enable_391), .CD(n14340), 
            .CK(clk_N_875), .Q(PWMdut_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i2 (.D(n2261[2]), .SP(clk_N_875_enable_391), .CD(n14336), 
            .CK(clk_N_875), .Q(PWMdut_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i1 (.D(n2261[1]), .SP(clk_N_875_enable_391), .CD(n14336), 
            .CK(clk_N_875), .Q(PWMdut_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i1.GSR = "DISABLED";
    FD1P3IX intgOut3_i28 (.D(intgOut0_28__N_1627[28]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i28.GSR = "ENABLED";
    FD1P3IX intgOut3_i27 (.D(intgOut0_28__N_1627[27]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i27.GSR = "ENABLED";
    FD1P3IX intgOut3_i26 (.D(intgOut0_28__N_1627[26]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i26.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i7 (.D0(n615[6]), .D1(addIn2_28__N_1569[6]), 
            .SD(n20384), .Z(addIn2_28__N_1440[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut3_i25 (.D(intgOut0_28__N_1627[25]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i25.GSR = "ENABLED";
    FD1P3IX intgOut3_i24 (.D(intgOut0_28__N_1627[24]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i24.GSR = "ENABLED";
    FD1P3IX intgOut3_i23 (.D(intgOut0_28__N_1627[23]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i23.GSR = "ENABLED";
    FD1P3IX intgOut3_i22 (.D(intgOut0_28__N_1627[22]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i22.GSR = "ENABLED";
    FD1P3IX intgOut3_i21 (.D(intgOut0_28__N_1627[21]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i21.GSR = "ENABLED";
    CCU2D sub_16_rep_4_add_2_13 (.A0(n4417), .B0(n11474), .C0(n5826), 
          .D0(n16073), .A1(n4416), .B1(n11474), .C1(n5828), .D1(n16073), 
          .CIN(n18674), .COUT(n18675), .S0(n4489), .S1(n4488));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_13.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_13.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_13.INJECT1_1 = "NO";
    FD1P3IX intgOut3_i20 (.D(intgOut0_28__N_1627[20]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i20.GSR = "ENABLED";
    FD1P3IX intgOut3_i19 (.D(intgOut0_28__N_1627[19]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i19.GSR = "ENABLED";
    FD1P3IX intgOut3_i18 (.D(intgOut0_28__N_1627[18]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i18.GSR = "ENABLED";
    FD1P3IX intgOut3_i17 (.D(intgOut0_28__N_1627[17]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i17.GSR = "ENABLED";
    FD1P3IX intgOut3_i16 (.D(intgOut0_28__N_1627[16]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i16.GSR = "ENABLED";
    FD1P3IX intgOut3_i15 (.D(intgOut0_28__N_1627[15]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i15.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i29 (.D0(n615[28]), .D1(addIn2_28__N_1569[28]), 
            .SD(n20384), .Z(addIn2_28__N_1440[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut3_i14 (.D(intgOut0_28__N_1627[14]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i14.GSR = "ENABLED";
    FD1P3IX intgOut3_i13 (.D(intgOut0_28__N_1627[13]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i13.GSR = "ENABLED";
    FD1P3IX intgOut3_i12 (.D(intgOut0_28__N_1627[12]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i12.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i8 (.D0(n615[7]), .D1(addIn2_28__N_1569[7]), 
            .SD(n20384), .Z(addIn2_28__N_1440[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut3_i11 (.D(intgOut0_28__N_1627[11]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i11.GSR = "ENABLED";
    FD1P3IX intgOut3_i10 (.D(intgOut0_28__N_1627[10]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i10.GSR = "ENABLED";
    FD1P3IX intgOut3_i9 (.D(intgOut0_28__N_1627[9]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i9.GSR = "ENABLED";
    FD1P3IX intgOut3_i8 (.D(intgOut0_28__N_1627[8]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i8.GSR = "ENABLED";
    CCU2D sub_16_rep_4_add_2_11 (.A0(n4419), .B0(n11474), .C0(n5822), 
          .D0(n16073), .A1(n4418), .B1(n11474), .C1(n5824), .D1(n16073), 
          .CIN(n18673), .COUT(n18674), .S0(n4491), .S1(n4490));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_11.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_11.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_11.INJECT1_1 = "NO";
    FD1P3IX intgOut3_i7 (.D(intgOut0_28__N_1627[7]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i7.GSR = "ENABLED";
    FD1P3IX intgOut3_i6 (.D(intgOut0_28__N_1627[6]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i6.GSR = "ENABLED";
    FD1P3IX intgOut3_i5 (.D(intgOut0_28__N_1627[5]), .SP(clk_N_875_enable_309), 
            .CD(n14313), .CK(clk_N_875), .Q(intgOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i5.GSR = "ENABLED";
    FD1P3IX intgOut2_i28 (.D(intgOut0_28__N_1627[28]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i28.GSR = "ENABLED";
    FD1P3IX intgOut2_i27 (.D(intgOut0_28__N_1627[27]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i27.GSR = "ENABLED";
    FD1P3IX intgOut2_i26 (.D(intgOut0_28__N_1627[26]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i26.GSR = "ENABLED";
    FD1P3IX intgOut2_i25 (.D(intgOut0_28__N_1627[25]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i25.GSR = "ENABLED";
    FD1P3IX intgOut2_i24 (.D(intgOut0_28__N_1627[24]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i24.GSR = "ENABLED";
    FD1P3IX intgOut2_i23 (.D(intgOut0_28__N_1627[23]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i23.GSR = "ENABLED";
    FD1P3IX intgOut2_i22 (.D(intgOut0_28__N_1627[22]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i22.GSR = "ENABLED";
    FD1P3IX intgOut2_i21 (.D(intgOut0_28__N_1627[21]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i21.GSR = "ENABLED";
    FD1P3IX intgOut2_i20 (.D(intgOut0_28__N_1627[20]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i20.GSR = "ENABLED";
    FD1P3IX intgOut2_i19 (.D(intgOut0_28__N_1627[19]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i19.GSR = "ENABLED";
    FD1P3IX intgOut2_i18 (.D(intgOut0_28__N_1627[18]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i18.GSR = "ENABLED";
    FD1P3IX intgOut2_i17 (.D(intgOut0_28__N_1627[17]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i17.GSR = "ENABLED";
    FD1P3IX intgOut2_i16 (.D(intgOut0_28__N_1627[16]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i16.GSR = "ENABLED";
    FD1P3IX intgOut2_i15 (.D(intgOut0_28__N_1627[15]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i15.GSR = "ENABLED";
    FD1P3IX intgOut2_i14 (.D(intgOut0_28__N_1627[14]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i14.GSR = "ENABLED";
    FD1P3IX intgOut2_i13 (.D(intgOut0_28__N_1627[13]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i13.GSR = "ENABLED";
    FD1P3IX intgOut2_i12 (.D(intgOut0_28__N_1627[12]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i12.GSR = "ENABLED";
    FD1P3IX intgOut2_i11 (.D(intgOut0_28__N_1627[11]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i11.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i9 (.D0(n615[8]), .D1(addIn2_28__N_1569[8]), 
            .SD(n20384), .Z(addIn2_28__N_1440[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut2_i10 (.D(intgOut0_28__N_1627[10]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i10.GSR = "ENABLED";
    FD1P3IX intgOut2_i9 (.D(intgOut0_28__N_1627[9]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i9.GSR = "ENABLED";
    FD1P3IX intgOut2_i8 (.D(intgOut0_28__N_1627[8]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i8.GSR = "ENABLED";
    FD1P3IX intgOut2_i7 (.D(intgOut0_28__N_1627[7]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i7.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i10 (.D0(n615[9]), .D1(addIn2_28__N_1569[9]), 
            .SD(n20384), .Z(addIn2_28__N_1440[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut2_i6 (.D(intgOut0_28__N_1627[6]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i6.GSR = "ENABLED";
    LUT4 i2_4_lut_else_3_lut_4_lut (.A(n22440), .B(ss[2]), .C(ss[3]), 
         .D(ss[0]), .Z(n22420)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam i2_4_lut_else_3_lut_4_lut.init = 16'hfffb;
    FD1P3IX intgOut2_i5 (.D(intgOut0_28__N_1627[5]), .SP(clk_N_875_enable_333), 
            .CD(n14289), .CK(clk_N_875), .Q(intgOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i5.GSR = "ENABLED";
    CCU2D sub_16_rep_4_add_2_9 (.A0(n4421), .B0(n11474), .C0(n5818), .D0(n16073), 
          .A1(n4420), .B1(n11474), .C1(n5820), .D1(n16073), .CIN(n18672), 
          .COUT(n18673), .S0(n4493), .S1(n4492));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_9.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_9.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_9.INJECT1_1 = "NO";
    FD1P3IX intgOut1_i28 (.D(intgOut0_28__N_1627[28]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i28.GSR = "ENABLED";
    FD1P3IX intgOut1_i27 (.D(intgOut0_28__N_1627[27]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i27.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_355_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n22433), 
         .D(n21729), .Z(n21668)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_355_3_lut_4_lut.init = 16'h0060;
    FD1P3IX intgOut1_i26 (.D(intgOut0_28__N_1627[26]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i26.GSR = "ENABLED";
    FD1P3IX intgOut1_i25 (.D(intgOut0_28__N_1627[25]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i25.GSR = "ENABLED";
    FD1P3IX intgOut1_i24 (.D(intgOut0_28__N_1627[24]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i24.GSR = "ENABLED";
    FD1P3IX intgOut1_i23 (.D(intgOut0_28__N_1627[23]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i23.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i11 (.D0(n615[10]), .D1(addIn2_28__N_1569[10]), 
            .SD(n20384), .Z(addIn2_28__N_1440[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_1_lut_rep_395 (.A(ss[0]), .Z(n21708)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut_rep_395.init = 16'h5555;
    FD1P3IX intgOut1_i22 (.D(intgOut0_28__N_1627[22]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i22.GSR = "ENABLED";
    FD1P3IX intgOut1_i21 (.D(intgOut0_28__N_1627[21]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i21.GSR = "ENABLED";
    FD1P3IX intgOut1_i20 (.D(intgOut0_28__N_1627[20]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i20.GSR = "ENABLED";
    LUT4 i13278_2_lut (.A(addOut[22]), .B(n22440), .Z(backOut3_28__N_1872[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13278_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_347_4_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(n21697), 
         .D(n22440), .Z(n21660)) /* synthesis lut_function=(!(A+(B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i1_2_lut_rep_347_4_lut_4_lut.init = 16'h0014;
    FD1P3IX intgOut1_i19 (.D(intgOut0_28__N_1627[19]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i19.GSR = "ENABLED";
    LUT4 i13102_2_lut_3_lut_3_lut_2_lut (.A(ss[0]), .B(n21674), .Z(multIn2[10])) /* synthesis lut_function=(A (B)) */ ;
    defparam i13102_2_lut_3_lut_3_lut_2_lut.init = 16'h8888;
    FD1P3IX intgOut1_i18 (.D(intgOut0_28__N_1627[18]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i18.GSR = "ENABLED";
    FD1P3IX intgOut1_i17 (.D(intgOut0_28__N_1627[17]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i17.GSR = "ENABLED";
    FD1P3IX intgOut1_i16 (.D(intgOut0_28__N_1627[16]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i16.GSR = "ENABLED";
    FD1P3IX intgOut1_i15 (.D(intgOut0_28__N_1627[15]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i15.GSR = "ENABLED";
    FD1P3IX intgOut1_i14 (.D(intgOut0_28__N_1627[14]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i14.GSR = "ENABLED";
    FD1P3IX intgOut1_i13 (.D(intgOut0_28__N_1627[13]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i13.GSR = "ENABLED";
    FD1P3IX intgOut1_i12 (.D(intgOut0_28__N_1627[12]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i12.GSR = "ENABLED";
    FD1P3IX intgOut1_i11 (.D(intgOut0_28__N_1627[11]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i11.GSR = "ENABLED";
    FD1P3IX intgOut1_i10 (.D(intgOut0_28__N_1627[10]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i10.GSR = "ENABLED";
    LUT4 i1_3_lut_adj_112 (.A(n1357[15]), .B(n2297[9]), .C(n30_adj_2327), 
         .Z(n19337)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[4] 376[11])
    defparam i1_3_lut_adj_112.init = 16'h8a8a;
    FD1P3IX intgOut1_i9 (.D(intgOut0_28__N_1627[9]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i9.GSR = "ENABLED";
    FD1P3IX intgOut1_i8 (.D(intgOut0_28__N_1627[8]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i8.GSR = "ENABLED";
    FD1P3IX intgOut1_i7 (.D(intgOut0_28__N_1627[7]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i7.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i12 (.D0(n615[11]), .D1(addIn2_28__N_1569[11]), 
            .SD(n20384), .Z(addIn2_28__N_1440[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i6 (.D(intgOut0_28__N_1627[6]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i6.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_113 (.A(n9_adj_2370), .B(n7_adj_2371), .C(n1357[10]), 
         .D(n1357[13]), .Z(n30_adj_2327)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_113.init = 16'h8000;
    FD1P3IX intgOut1_i5 (.D(intgOut0_28__N_1627[5]), .SP(clk_N_875_enable_392), 
            .CD(n14265), .CK(clk_N_875), .Q(intgOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i5.GSR = "ENABLED";
    FD1P3IX intgOut1_i4 (.D(addOut[4]), .SP(clk_N_875_enable_392), .CD(n14260), 
            .CK(clk_N_875), .Q(intgOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i4.GSR = "ENABLED";
    FD1P3IX intgOut1_i3 (.D(addOut[3]), .SP(clk_N_875_enable_392), .CD(n14260), 
            .CK(clk_N_875), .Q(intgOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i3.GSR = "ENABLED";
    FD1P3IX intgOut1_i2 (.D(addOut[2]), .SP(clk_N_875_enable_392), .CD(n14260), 
            .CK(clk_N_875), .Q(intgOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i2.GSR = "ENABLED";
    FD1P3IX intgOut1_i1 (.D(addOut[1]), .SP(clk_N_875_enable_392), .CD(n14260), 
            .CK(clk_N_875), .Q(intgOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i1.GSR = "ENABLED";
    FD1P3IX intgOut0_i28 (.D(intgOut0_28__N_1627[28]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i28.GSR = "ENABLED";
    FD1P3IX intgOut0_i27 (.D(intgOut0_28__N_1627[27]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i27.GSR = "ENABLED";
    PFUMX i17636 (.BLUT(n21515), .ALUT(n21677), .C0(n22440), .Z(clk_N_875_enable_136));
    FD1P3IX intgOut0_i26 (.D(intgOut0_28__N_1627[26]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i26.GSR = "ENABLED";
    FD1P3IX intgOut0_i25 (.D(intgOut0_28__N_1627[25]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i25.GSR = "ENABLED";
    FD1P3IX intgOut0_i24 (.D(intgOut0_28__N_1627[24]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i24.GSR = "ENABLED";
    FD1P3IX intgOut0_i23 (.D(intgOut0_28__N_1627[23]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i23.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i13 (.D0(n615[12]), .D1(addIn2_28__N_1569[12]), 
            .SD(n20384), .Z(addIn2_28__N_1440[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i22 (.D(intgOut0_28__N_1627[22]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i22.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i14 (.D0(n615[13]), .D1(addIn2_28__N_1569[13]), 
            .SD(n20384), .Z(addIn2_28__N_1440[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i15 (.D0(n615[14]), .D1(addIn2_28__N_1569[14]), 
            .SD(n20384), .Z(addIn2_28__N_1440[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i21 (.D(intgOut0_28__N_1627[21]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i21.GSR = "ENABLED";
    FD1P3IX intgOut0_i20 (.D(intgOut0_28__N_1627[20]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i20.GSR = "ENABLED";
    FD1P3IX intgOut0_i19 (.D(intgOut0_28__N_1627[19]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i19.GSR = "ENABLED";
    FD1P3IX intgOut0_i18 (.D(intgOut0_28__N_1627[18]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i18.GSR = "ENABLED";
    FD1P3IX intgOut0_i17 (.D(intgOut0_28__N_1627[17]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i17.GSR = "ENABLED";
    FD1P3IX intgOut0_i16 (.D(intgOut0_28__N_1627[16]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i16.GSR = "ENABLED";
    FD1P3IX intgOut0_i15 (.D(intgOut0_28__N_1627[15]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i15.GSR = "ENABLED";
    FD1P3IX intgOut0_i14 (.D(intgOut0_28__N_1627[14]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i14.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i16 (.D0(n615[15]), .D1(addIn2_28__N_1569[15]), 
            .SD(n20384), .Z(addIn2_28__N_1440[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i13 (.D(intgOut0_28__N_1627[13]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i13.GSR = "ENABLED";
    LUT4 i3_2_lut_adj_114 (.A(n1357[14]), .B(n1357[12]), .Z(n9_adj_2370)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_114.init = 16'h8888;
    FD1P3IX intgOut0_i12 (.D(intgOut0_28__N_1627[12]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i12.GSR = "ENABLED";
    FD1P3IX intgOut0_i11 (.D(intgOut0_28__N_1627[11]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i11.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i17 (.D0(n615[16]), .D1(addIn2_28__N_1569[16]), 
            .SD(n20384), .Z(addIn2_28__N_1440[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i10 (.D(intgOut0_28__N_1627[10]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i10.GSR = "ENABLED";
    FD1P3IX intgOut0_i9 (.D(intgOut0_28__N_1627[9]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i9.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i18 (.D0(n615[17]), .D1(addIn2_28__N_1569[17]), 
            .SD(n20384), .Z(addIn2_28__N_1440[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i8 (.D(intgOut0_28__N_1627[8]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i8.GSR = "ENABLED";
    FD1P3IX intgOut0_i7 (.D(intgOut0_28__N_1627[7]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i7.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i19 (.D0(n615[18]), .D1(addIn2_28__N_1569[18]), 
            .SD(n20384), .Z(addIn2_28__N_1440[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i6 (.D(intgOut0_28__N_1627[6]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i6.GSR = "ENABLED";
    FD1P3IX intgOut0_i5 (.D(intgOut0_28__N_1627[5]), .SP(clk_N_875_enable_389), 
            .CD(n14237), .CK(clk_N_875), .Q(intgOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i5.GSR = "ENABLED";
    FD1P3IX intgOut0_i4 (.D(addOut[4]), .SP(clk_N_875_enable_389), .CD(n14232), 
            .CK(clk_N_875), .Q(intgOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i4.GSR = "ENABLED";
    FD1P3IX intgOut0_i3 (.D(addOut[3]), .SP(clk_N_875_enable_389), .CD(n14232), 
            .CK(clk_N_875), .Q(intgOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i3.GSR = "ENABLED";
    FD1P3IX intgOut0_i2 (.D(addOut[2]), .SP(clk_N_875_enable_389), .CD(n14232), 
            .CK(clk_N_875), .Q(intgOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i2.GSR = "ENABLED";
    FD1P3IX intgOut0_i1 (.D(addOut[1]), .SP(clk_N_875_enable_389), .CD(n14232), 
            .CK(clk_N_875), .Q(intgOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i1.GSR = "ENABLED";
    L6MUX21 addIn2_28__I_29_i20 (.D0(n615[19]), .D1(addIn2_28__N_1569[19]), 
            .SD(n20384), .Z(addIn2_28__N_1440[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_4_lut_adj_115 (.A(n1357[11]), .B(n1357[9]), .C(n10_adj_2372), 
         .D(n1357[7]), .Z(n7_adj_2371)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_115.init = 16'haaa8;
    L6MUX21 addIn2_28__I_29_i21 (.D0(n615[20]), .D1(addIn2_28__N_1569[20]), 
            .SD(n20384), .Z(addIn2_28__N_1440[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i22 (.D0(n615[21]), .D1(addIn2_28__N_1569[21]), 
            .SD(n20384), .Z(addIn2_28__N_1440[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i23 (.D0(n615[22]), .D1(addIn2_28__N_1569[22]), 
            .SD(n20384), .Z(addIn2_28__N_1440[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1S3IX ss_i2_rep_424 (.D(n14), .CK(clk_N_875), .CD(ss[4]), .Q(n22433));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i2_rep_424.GSR = "ENABLED";
    LUT4 i13498_2_lut (.A(addOut[21]), .B(n22440), .Z(Out2_28__N_1145[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13498_2_lut.init = 16'h2222;
    LUT4 i4_4_lut_adj_116 (.A(n1357[6]), .B(n8_adj_2373), .C(n1357[4]), 
         .D(n4_adj_2374), .Z(n10_adj_2372)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_116.init = 16'hfeee;
    L6MUX21 addIn2_28__I_29_i2 (.D0(n615[1]), .D1(addIn2_28__N_1569[1]), 
            .SD(n20384), .Z(addIn2_28__N_1440[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D sub_16_rep_4_add_2_7 (.A0(n4423), .B0(n11474), .C0(n5814), .D0(n16073), 
          .A1(n4422), .B1(n11474), .C1(n5816), .D1(n16073), .CIN(n18671), 
          .COUT(n18672), .S0(n4495), .S1(n4494));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_7.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_7.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_7.INJECT1_1 = "NO";
    LUT4 i2_2_lut_adj_117 (.A(n1357[5]), .B(n1357[8]), .Z(n8_adj_2373)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_117.init = 16'heeee;
    L6MUX21 addIn2_28__I_29_i24 (.D0(n615[23]), .D1(addIn2_28__N_1569[23]), 
            .SD(n20384), .Z(addIn2_28__N_1440[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_4_lut_adj_118 (.A(n1357[3]), .B(n1357[2]), .C(n1357[1]), .D(n1357[0]), 
         .Z(n4_adj_2374)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_118.init = 16'haaa8;
    L6MUX21 addIn2_28__I_29_i3 (.D0(n615[2]), .D1(addIn2_28__N_1569[2]), 
            .SD(n20384), .Z(addIn2_28__N_1440[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i1 (.D0(n615[0]), .D1(addIn2_28__N_1569[0]), 
            .SD(n20384), .Z(addIn2_28__N_1440[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i13 (.BLUT(n367[12]), .ALUT(subIn2_24__N_1348[12]), 
          .C0(n20645), .Z(n4416)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i10 (.BLUT(n367[9]), .ALUT(subIn2_24__N_1348[9]), 
          .C0(n20645), .Z(n4419)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_3_lut_adj_119 (.A(n1357[15]), .B(n2297[8]), .C(n30_adj_2327), 
         .Z(n19331)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[4] 376[11])
    defparam i1_3_lut_adj_119.init = 16'h8a8a;
    PFUMX subIn2_24__I_0_rep_1_i9 (.BLUT(n367[8]), .ALUT(subIn2_24__N_1348[8]), 
          .C0(n20645), .Z(n4420)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i8 (.BLUT(n367[7]), .ALUT(subIn2_24__N_1348[7]), 
          .C0(n20645), .Z(n4421)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i4 (.BLUT(n367[3]), .ALUT(subIn2_24__N_1348[3]), 
          .C0(n20645), .Z(n4425)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i20 (.BLUT(subIn2_24__N_1534[19]), .ALUT(subIn2_24__N_1348[19]), 
          .C0(n20659), .Z(n4409)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_3_lut_adj_120 (.A(n1357[15]), .B(n2297[7]), .C(n30_adj_2327), 
         .Z(n19325)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[4] 376[11])
    defparam i1_3_lut_adj_120.init = 16'h8a8a;
    PFUMX subIn2_24__I_0_rep_1_i19 (.BLUT(subIn2_24__N_1534[18]), .ALUT(subIn2_24__N_1348[18]), 
          .C0(n20659), .Z(n4410)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13274_2_lut (.A(addOut[20]), .B(n22440), .Z(backOut3_28__N_1872[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13274_2_lut.init = 16'h2222;
    PFUMX subIn2_24__I_0_rep_1_i18 (.BLUT(subIn2_24__N_1534[17]), .ALUT(subIn2_24__N_1348[17]), 
          .C0(n20659), .Z(n4411)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_189_i19_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[18]), 
         .Z(intgOut0_28__N_1627[18])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i19_3_lut_3_lut.init = 16'hbaba;
    PFUMX subIn2_24__I_0_rep_1_i17 (.BLUT(subIn2_24__N_1534[16]), .ALUT(subIn2_24__N_1348[16]), 
          .C0(n20659), .Z(n4412)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_1253_i21_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[20]), 
         .D(speed_set_m4[20]), .Z(n2593[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1253_i3_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[2]), 
         .D(speed_set_m4[2]), .Z(n2593[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_adj_121 (.A(n1357[15]), .B(n2297[6]), .C(n30_adj_2327), 
         .Z(n1539[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_121.init = 16'h8a8a;
    PFUMX subIn2_24__I_0_rep_1_i16 (.BLUT(subIn2_24__N_1534[15]), .ALUT(subIn2_24__N_1348[15]), 
          .C0(n20659), .Z(n4413)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_189_i18_3_lut_3_lut (.A(n1065), .B(n3844), .C(addOut[17]), 
         .Z(intgOut0_28__N_1627[17])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i18_3_lut_3_lut.init = 16'hbaba;
    LUT4 i1_3_lut_adj_122 (.A(n1357[15]), .B(n2297[5]), .C(n30_adj_2327), 
         .Z(n1539[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_122.init = 16'h8a8a;
    LUT4 mux_1253_i7_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[6]), 
         .D(speed_set_m4[6]), .Z(n2593[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1253_i2_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[1]), 
         .D(speed_set_m4[1]), .Z(n2593[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i2_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_rep_315_3_lut (.A(n1065), .B(n3844), .C(n22440), .Z(n21628)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_315_3_lut.init = 16'hfefe;
    PFUMX subIn2_24__I_0_rep_1_i15 (.BLUT(subIn2_24__N_1534[14]), .ALUT(subIn2_24__N_1348[14]), 
          .C0(n20659), .Z(n4414)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_3_lut_adj_123 (.A(n1336[15]), .B(n2285[9]), .C(n9_adj_2375), 
         .Z(n1495[9])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_123.init = 16'h8a8a;
    PFUMX subIn2_24__I_0_rep_1_i14 (.BLUT(subIn2_24__N_1534[13]), .ALUT(subIn2_24__N_1348[13]), 
          .C0(n20659), .Z(n4415)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_215_17 (.A0(Out1[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18436), 
          .S0(n1315[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_17.INIT0 = 16'h5aaa;
    defparam add_215_17.INIT1 = 16'h0000;
    defparam add_215_17.INJECT1_0 = "NO";
    defparam add_215_17.INJECT1_1 = "NO";
    PFUMX subIn2_24__I_0_rep_1_i12 (.BLUT(subIn2_24__N_1534[11]), .ALUT(subIn2_24__N_1348[11]), 
          .C0(n20659), .Z(n4417)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i5_4_lut_adj_124 (.A(n9_adj_2376), .B(n1336[10]), .C(n8_adj_2377), 
         .D(n1336[11]), .Z(n9_adj_2375)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_124.init = 16'h8000;
    PFUMX subIn2_24__I_0_rep_1_i11 (.BLUT(subIn2_24__N_1534[10]), .ALUT(subIn2_24__N_1348[10]), 
          .C0(n20659), .Z(n4418)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i7 (.BLUT(subIn2_24__N_1534[6]), .ALUT(subIn2_24__N_1348[6]), 
          .C0(n20659), .Z(n4422)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13030_2_lut_rep_408 (.A(ss[0]), .B(ss[1]), .Z(n21721)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13030_2_lut_rep_408.init = 16'h8888;
    PFUMX subIn2_24__I_0_rep_1_i6 (.BLUT(subIn2_24__N_1534[5]), .ALUT(subIn2_24__N_1348[5]), 
          .C0(n20659), .Z(n4423)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13495_2_lut (.A(addOut[18]), .B(n22440), .Z(Out2_28__N_1145[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13495_2_lut.init = 16'h2222;
    PFUMX subIn2_24__I_0_rep_1_i5 (.BLUT(subIn2_24__N_1534[4]), .ALUT(subIn2_24__N_1348[4]), 
          .C0(n20659), .Z(n4424)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i3 (.BLUT(subIn2_24__N_1534[2]), .ALUT(subIn2_24__N_1348[2]), 
          .C0(n20659), .Z(n4426)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i2 (.BLUT(subIn2_24__N_1534[1]), .ALUT(subIn2_24__N_1348[1]), 
          .C0(n20659), .Z(n4427)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i1 (.BLUT(subIn2_24__N_1534[0]), .ALUT(subIn2_24__N_1348[0]), 
          .C0(n20659), .Z(n4428)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i9 (.BLUT(n555[8]), .ALUT(n675[8]), .C0(n20372), .Z(addIn2_28__N_1569[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i10 (.BLUT(n555[9]), .ALUT(n675[9]), .C0(n20372), .Z(addIn2_28__N_1569[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i11 (.BLUT(n555[10]), .ALUT(n675[10]), .C0(n20372), 
          .Z(addIn2_28__N_1569[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_1253_i9_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[8]), 
         .D(speed_set_m4[8]), .Z(n2593[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i9_3_lut_4_lut.init = 16'hfe10;
    PFUMX mux_140_i12 (.BLUT(n555[11]), .ALUT(n675[11]), .C0(n20372), 
          .Z(addIn2_28__N_1569[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i13 (.BLUT(n555[12]), .ALUT(n675[12]), .C0(n20372), 
          .Z(addIn2_28__N_1569[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i3_2_lut_adj_125 (.A(n1336[14]), .B(n1336[13]), .Z(n9_adj_2376)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_125.init = 16'h8888;
    LUT4 i2_4_lut_adj_126 (.A(n1336[9]), .B(n1336[12]), .C(n10_adj_2378), 
         .D(n1336[7]), .Z(n8_adj_2377)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_126.init = 16'hccc8;
    LUT4 i4_4_lut_adj_127 (.A(n1336[6]), .B(n8_adj_2379), .C(n1336[4]), 
         .D(n4_adj_2380), .Z(n10_adj_2378)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_127.init = 16'hfeee;
    LUT4 i2_2_lut_adj_128 (.A(n1336[5]), .B(n1336[8]), .Z(n8_adj_2379)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_128.init = 16'heeee;
    PFUMX mux_140_i14 (.BLUT(n555[13]), .ALUT(n675[13]), .C0(n20372), 
          .Z(addIn2_28__N_1569[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_4_lut_adj_129 (.A(n1336[3]), .B(n1336[2]), .C(n1336[1]), .D(n1336[0]), 
         .Z(n4_adj_2380)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_129.init = 16'haaa8;
    PFUMX mux_140_i15 (.BLUT(n555[14]), .ALUT(n675[14]), .C0(n20372), 
          .Z(addIn2_28__N_1569[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i16 (.BLUT(n555[15]), .ALUT(n675[15]), .C0(n20372), 
          .Z(addIn2_28__N_1569[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i17 (.BLUT(n555[16]), .ALUT(n675[16]), .C0(n20372), 
          .Z(addIn2_28__N_1569[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i18 (.BLUT(n555[17]), .ALUT(n675[17]), .C0(n20372), 
          .Z(addIn2_28__N_1569[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i19 (.BLUT(n555[18]), .ALUT(n675[18]), .C0(n20372), 
          .Z(addIn2_28__N_1569[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i20 (.BLUT(n555[19]), .ALUT(n675[19]), .C0(n20372), 
          .Z(addIn2_28__N_1569[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i21 (.BLUT(n555[20]), .ALUT(n675[20]), .C0(n20372), 
          .Z(addIn2_28__N_1569[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_3_lut_adj_130 (.A(n1336[15]), .B(n2285[8]), .C(n9_adj_2375), 
         .Z(n1495[8])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_130.init = 16'h8a8a;
    LUT4 equal_110_i9_2_lut_rep_353_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n22425), 
         .D(ss[3]), .Z(n21666)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam equal_110_i9_2_lut_rep_353_3_lut_4_lut.init = 16'hf7ff;
    PFUMX mux_140_i22 (.BLUT(n555[21]), .ALUT(n675[21]), .C0(n20372), 
          .Z(addIn2_28__N_1569[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13582_2_lut_rep_319_3_lut (.A(n22411), .B(n22440), .C(n56), 
         .Z(n21632)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i13582_2_lut_rep_319_3_lut.init = 16'hfefe;
    PFUMX mux_140_i23 (.BLUT(n555[22]), .ALUT(n675[22]), .C0(n20372), 
          .Z(addIn2_28__N_1569[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i7928_2_lut_3_lut (.A(ss[0]), .B(ss[1]), .C(ss[2]), .Z(n14)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i7928_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_3_lut_adj_131 (.A(n1336[15]), .B(n2285[7]), .C(n9_adj_2375), 
         .Z(n1495[7])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_131.init = 16'h8a8a;
    LUT4 i1_3_lut_adj_132 (.A(n1336[15]), .B(n2285[6]), .C(n9_adj_2375), 
         .Z(n1495[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_132.init = 16'h8a8a;
    LUT4 mux_1253_i16_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[15]), 
         .D(speed_set_m4[15]), .Z(n2593[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3_2_lut_3_lut_4_lut (.A(n22411), .B(n22440), .C(subIn1_24__N_1342), 
         .D(n56), .Z(n8_adj_2369)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i3_2_lut_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i1_3_lut_adj_133 (.A(n1315[15]), .B(n2273[5]), .C(n30), .Z(n1451[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_133.init = 16'h8a8a;
    LUT4 mux_138_i9_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[8]), 
         .D(intgOut2[8]), .Z(n645[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i9_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_4_lut_adj_134 (.A(n16469), .B(n16127), .C(n21677), .D(n22440), 
         .Z(clk_N_875_enable_333)) /* synthesis lut_function=((B (C (D))+!B (C+!(D)))+!A) */ ;
    defparam i1_4_lut_adj_134.init = 16'hf577;
    LUT4 i1855_2_lut_rep_418 (.A(ss[0]), .B(ss[1]), .Z(n22419)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1855_2_lut_rep_418.init = 16'h6666;
    LUT4 i2_3_lut_rep_335_4_lut_then_3_lut (.A(ss[3]), .B(n22425), .C(ss[1]), 
         .Z(n22427)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(174[9:17])
    defparam i2_3_lut_rep_335_4_lut_then_3_lut.init = 16'hdfdf;
    LUT4 i16724_2_lut_rep_421 (.A(n22433), .B(n22440), .Z(n22425)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16724_2_lut_rep_421.init = 16'heeee;
    LUT4 i1_3_lut_adj_135 (.A(n1336[15]), .B(n2285[5]), .C(n9_adj_2375), 
         .Z(n1495[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_135.init = 16'h8a8a;
    LUT4 n15590_bdd_4_lut_rep_419 (.A(n21729), .B(ss[0]), .C(n22433), 
         .D(ss[1]), .Z(n22423)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam n15590_bdd_4_lut_rep_419.init = 16'h0410;
    LUT4 i2_4_lut_then_3_lut_4_lut (.A(ss[2]), .B(n22440), .C(ss[3]), 
         .D(ss[0]), .Z(n22421)) /* synthesis lut_function=(A+(B+(C (D)+!C !(D)))) */ ;
    defparam i2_4_lut_then_3_lut_4_lut.init = 16'hfeef;
    LUT4 i1_4_lut_adj_136 (.A(n3708), .B(n35_adj_2381), .C(n40_adj_2382), 
         .D(n36_adj_2383), .Z(n4_adj_2338)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_136.init = 16'haaa8;
    PFUMX mux_140_i24 (.BLUT(n555[23]), .ALUT(n675[23]), .C0(n20372), 
          .Z(addIn2_28__N_1569[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i25 (.BLUT(n555[24]), .ALUT(n675[24]), .C0(n20372), 
          .Z(addIn2_28__N_1569[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i2 (.BLUT(n555[1]), .ALUT(n675[1]), .C0(n20372), .Z(addIn2_28__N_1569[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i26 (.BLUT(n555[25]), .ALUT(n675[25]), .C0(n20372), 
          .Z(addIn2_28__N_1569[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i3 (.BLUT(n555[2]), .ALUT(n675[2]), .C0(n20372), .Z(addIn2_28__N_1569[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i27 (.BLUT(n555[26]), .ALUT(n675[26]), .C0(n20372), 
          .Z(addIn2_28__N_1569[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_3_lut_adj_137 (.A(n1315[15]), .B(n2273[3]), .C(n30), .Z(n1451[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_137.init = 16'h8a8a;
    LUT4 i1_4_lut_then_4_lut (.A(n22440), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21737)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0040;
    FD1P3IX dutyout_m4_i0_i0 (.D(n2297[0]), .SP(clk_N_875_enable_391), .CD(n14363), 
            .CK(clk_N_875), .Q(PWMdut_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i0.GSR = "DISABLED";
    LUT4 i1_4_lut_else_4_lut (.A(n22440), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21736)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0100;
    PFUMX mux_140_i4 (.BLUT(n555[3]), .ALUT(n675[3]), .C0(n20372), .Z(addIn2_28__N_1569[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_1253_i10_3_lut_4_lut (.A(n15564), .B(n49), .C(speed_set_m3[9]), 
         .D(speed_set_m4[9]), .Z(n2593[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1253_i10_3_lut_4_lut.init = 16'hfe10;
    PFUMX mux_140_i28 (.BLUT(n555[27]), .ALUT(n675[27]), .C0(n20372), 
          .Z(addIn2_28__N_1569[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i5 (.BLUT(n555[4]), .ALUT(n675[4]), .C0(n20372), .Z(addIn2_28__N_1569[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX dutyout_m3_i0_i0 (.D(n2285[0]), .SP(clk_N_875_enable_391), .CD(n14354), 
            .CK(clk_N_875), .Q(PWMdut_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i0.GSR = "DISABLED";
    PFUMX mux_140_i29 (.BLUT(n555[28]), .ALUT(n675[28]), .C0(n20372), 
          .Z(addIn2_28__N_1569[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i14_4_lut_adj_138 (.A(speed_set_m3[13]), .B(speed_set_m3[1]), .C(speed_set_m3[12]), 
         .D(speed_set_m3[2]), .Z(n35_adj_2381)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_138.init = 16'hfffe;
    LUT4 i19_4_lut_adj_139 (.A(speed_set_m3[15]), .B(n38_adj_2384), .C(n32_adj_2385), 
         .D(speed_set_m3[10]), .Z(n40_adj_2382)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_139.init = 16'hfffe;
    LUT4 i15_4_lut_adj_140 (.A(speed_set_m3[0]), .B(speed_set_m3[7]), .C(speed_set_m3[17]), 
         .D(speed_set_m3[11]), .Z(n36_adj_2383)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_140.init = 16'hfffe;
    FD1P3IX intgOut1_i0 (.D(addOut[0]), .SP(clk_N_875_enable_392), .CD(n14260), 
            .CK(clk_N_875), .Q(intgOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i0.GSR = "ENABLED";
    LUT4 i17_4_lut_adj_141 (.A(speed_set_m3[8]), .B(n34_adj_2329), .C(n24_adj_2330), 
         .D(speed_set_m3[16]), .Z(n38_adj_2384)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_141.init = 16'hfffe;
    PFUMX mux_140_i6 (.BLUT(n555[5]), .ALUT(n675[5]), .C0(n20372), .Z(addIn2_28__N_1569[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13492_2_lut (.A(addOut[17]), .B(n22440), .Z(Out2_28__N_1145[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13492_2_lut.init = 16'h2222;
    PFUMX mux_140_i7 (.BLUT(n555[6]), .ALUT(n675[6]), .C0(n20372), .Z(addIn2_28__N_1569[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13487_2_lut (.A(addOut[16]), .B(n22440), .Z(Out2_28__N_1145[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13487_2_lut.init = 16'h2222;
    PFUMX mux_140_i8 (.BLUT(n555[7]), .ALUT(n675[7]), .C0(n20372), .Z(addIn2_28__N_1569[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i11769_4_lut (.A(clk_N_875_enable_391), .B(n1336[15]), .C(n9_adj_2375), 
         .D(n18943), .Z(n14354)) /* synthesis lut_function=(A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11769_4_lut.init = 16'haa2a;
    LUT4 i13484_2_lut (.A(addOut[15]), .B(n22440), .Z(Out2_28__N_1145[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13484_2_lut.init = 16'h2222;
    LUT4 n22411_bdd_2_lut_rep_417 (.A(n22411), .B(n22440), .Z(n22418)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n22411_bdd_2_lut_rep_417.init = 16'heeee;
    LUT4 i1_2_lut_rep_368_3_lut (.A(n22440), .B(ss[2]), .C(ss[3]), .Z(n21681)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam i1_2_lut_rep_368_3_lut.init = 16'hbfbf;
    LUT4 i13266_2_lut (.A(addOut[14]), .B(n22440), .Z(backOut3_28__N_1872[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13266_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_adj_142 (.A(n1336[15]), .B(n2285[3]), .C(n9_adj_2375), 
         .Z(n1495[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_142.init = 16'h8a8a;
    LUT4 i11_3_lut_adj_143 (.A(speed_set_m3[6]), .B(speed_set_m3[3]), .C(speed_set_m3[14]), 
         .Z(n32_adj_2385)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_143.init = 16'hfefe;
    LUT4 i13265_2_lut (.A(addOut[13]), .B(n22440), .Z(backOut3_28__N_1872[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13265_2_lut.init = 16'h2222;
    LUT4 equal_114_i9_2_lut_rep_346_3_lut_4_lut (.A(n22440), .B(ss[2]), 
         .C(n6), .D(ss[3]), .Z(n21659)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam equal_114_i9_2_lut_rep_346_3_lut_4_lut.init = 16'hfbff;
    LUT4 i1_3_lut_adj_144 (.A(n1315[15]), .B(n2273[9]), .C(n30), .Z(n19319)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[4] 360[11])
    defparam i1_3_lut_adj_144.init = 16'h8a8a;
    PFUMX mux_140_i1 (.BLUT(n555[0]), .ALUT(n675[0]), .C0(n20372), .Z(addIn2_28__N_1569[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13475_2_lut (.A(addOut[12]), .B(n22440), .Z(Out2_28__N_1145[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13475_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_adj_145 (.A(n1315[15]), .B(n2273[8]), .C(n30), .Z(n19313)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[4] 360[11])
    defparam i1_3_lut_adj_145.init = 16'h8a8a;
    PFUMX mux_137_i2 (.BLUT(n585[1]), .ALUT(intgOut3[1]), .C0(n21646), 
          .Z(n615[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13474_2_lut (.A(addOut[11]), .B(n22440), .Z(Out2_28__N_1145[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13474_2_lut.init = 16'h2222;
    PFUMX mux_137_i3 (.BLUT(n585[2]), .ALUT(intgOut3[2]), .C0(n21646), 
          .Z(n615[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i4 (.BLUT(n585[3]), .ALUT(intgOut3[3]), .C0(n21646), 
          .Z(n615[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i5 (.BLUT(n585[4]), .ALUT(intgOut3[4]), .C0(n21646), 
          .Z(n615[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 equal_133_i9_2_lut_3_lut_4_lut (.A(n22440), .B(n22433), .C(n21723), 
         .D(ss[3]), .Z(n9_adj_2331)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam equal_133_i9_2_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 i1_3_lut_adj_146 (.A(n1315[15]), .B(n2273[7]), .C(n30), .Z(n19307)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[4] 360[11])
    defparam i1_3_lut_adj_146.init = 16'h8a8a;
    PFUMX mux_137_i6 (.BLUT(n585[5]), .ALUT(intgOut3[5]), .C0(n21646), 
          .Z(n615[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i7 (.BLUT(n585[6]), .ALUT(intgOut3[6]), .C0(n21646), 
          .Z(n615[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i8 (.BLUT(n585[7]), .ALUT(intgOut3[7]), .C0(n21646), 
          .Z(n615[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i9 (.BLUT(n585[8]), .ALUT(intgOut3[8]), .C0(n21646), 
          .Z(n615[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i10 (.BLUT(n585[9]), .ALUT(intgOut3[9]), .C0(n21646), 
          .Z(n615[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i11 (.BLUT(n585[10]), .ALUT(intgOut3[10]), .C0(n21646), 
          .Z(n615[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 ss_4__I_0_351_i6_2_lut_rep_410 (.A(ss[0]), .B(ss[1]), .Z(n21723)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(164[29:36])
    defparam ss_4__I_0_351_i6_2_lut_rep_410.init = 16'hbbbb;
    PFUMX mux_137_i12 (.BLUT(n585[11]), .ALUT(intgOut3[11]), .C0(n21646), 
          .Z(n615[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_215_15 (.A0(Out1[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18435), 
          .COUT(n18436), .S0(n1315[13]), .S1(n1315[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_15.INIT0 = 16'h5aaa;
    defparam add_215_15.INIT1 = 16'h5aaa;
    defparam add_215_15.INJECT1_0 = "NO";
    defparam add_215_15.INJECT1_1 = "NO";
    PFUMX mux_137_i13 (.BLUT(n585[12]), .ALUT(intgOut3[12]), .C0(n21646), 
          .Z(n615[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13471_2_lut (.A(addOut[10]), .B(n22440), .Z(Out2_28__N_1145[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13471_2_lut.init = 16'h2222;
    PFUMX mux_137_i14 (.BLUT(n585[13]), .ALUT(intgOut3[13]), .C0(n21646), 
          .Z(n615[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_138_i10_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[9]), 
         .D(intgOut2[9]), .Z(n645[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i10_3_lut_4_lut.init = 16'hfe10;
    PFUMX mux_137_i15 (.BLUT(n585[14]), .ALUT(intgOut3[14]), .C0(n21646), 
          .Z(n615[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_138_i18_3_lut_4_lut (.A(n6), .B(n22424), .C(intgOut1[17]), 
         .D(intgOut2[17]), .Z(n645[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i18_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13255_2_lut (.A(addOut[9]), .B(n22440), .Z(backOut3_28__N_1872[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13255_2_lut.init = 16'h2222;
    PFUMX mux_137_i16 (.BLUT(n585[15]), .ALUT(intgOut3[15]), .C0(n21646), 
          .Z(n615[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i17 (.BLUT(n585[16]), .ALUT(intgOut3[16]), .C0(n21646), 
          .Z(n615[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i18 (.BLUT(n585[17]), .ALUT(intgOut3[17]), .C0(n21646), 
          .Z(n615[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i19 (.BLUT(n585[18]), .ALUT(intgOut3[18]), .C0(n21646), 
          .Z(n615[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i20 (.BLUT(n585[19]), .ALUT(intgOut3[19]), .C0(n21646), 
          .Z(n615[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i21 (.BLUT(n585[20]), .ALUT(intgOut3[20]), .C0(n21646), 
          .Z(n615[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D sub_16_rep_4_add_2_5 (.A0(n4425), .B0(n11474), .C0(n5810), .D0(n16073), 
          .A1(n4424), .B1(n11474), .C1(n5812), .D1(n16073), .CIN(n18670), 
          .COUT(n18671), .S0(n4497), .S1(n4496));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_5.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_5.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_3 (.A0(n4427), .B0(n11474), .C0(n5806), .D0(n16073), 
          .A1(n4426), .B1(n11474), .C1(n5808), .D1(n16073), .CIN(n18669), 
          .COUT(n18670), .S0(n4499), .S1(n4498));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_3.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_3.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n4428), .B1(n11474), .C1(n5519), .D1(n16073), 
          .COUT(n18669), .S1(n4500));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_1.INIT0 = 16'h0000;
    defparam sub_16_rep_4_add_2_1.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_1.INJECT1_1 = "NO";
    CCU2D add_211_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[13]), .B1(n18945), .C1(n18946), .D1(Out0[28]), .COUT(n18421), 
          .S1(n1294[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_1.INIT0 = 16'hF000;
    defparam add_211_1.INIT1 = 16'h56aa;
    defparam add_211_1.INJECT1_0 = "NO";
    defparam add_211_1.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_23 (.A0(n2353[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18667), .S0(n4454), .S1(n4453));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_23.INIT0 = 16'h5555;
    defparam sub_16_rep_3_add_2_23.INIT1 = 16'h5555;
    defparam sub_16_rep_3_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_23.INJECT1_1 = "NO";
    CCU2D add_215_13 (.A0(Out1[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18434), 
          .COUT(n18435), .S0(n1315[11]), .S1(n1315[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_13.INIT0 = 16'h5aaa;
    defparam add_215_13.INIT1 = 16'h5aaa;
    defparam add_215_13.INJECT1_0 = "NO";
    defparam add_215_13.INJECT1_1 = "NO";
    PFUMX mux_137_i22 (.BLUT(n585[21]), .ALUT(intgOut3[21]), .C0(n21646), 
          .Z(n615[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_1188_23 (.A0(n5450), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18420), 
          .S0(n2353[21]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_23.INIT0 = 16'hf555;
    defparam add_1188_23.INIT1 = 16'h0000;
    defparam add_1188_23.INJECT1_0 = "NO";
    defparam add_1188_23.INJECT1_1 = "NO";
    PFUMX mux_137_i1 (.BLUT(n585[0]), .ALUT(intgOut3[0]), .C0(n21646), 
          .Z(n615[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_1188_21 (.A0(n5448), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5450), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18419), 
          .COUT(n18420), .S0(n2353[19]), .S1(n2353[20]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_21.INIT0 = 16'hf555;
    defparam add_1188_21.INIT1 = 16'hf555;
    defparam add_1188_21.INJECT1_0 = "NO";
    defparam add_1188_21.INJECT1_1 = "NO";
    CCU2D add_215_11 (.A0(Out1[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18433), 
          .COUT(n18434), .S0(n1315[9]), .S1(n1315[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_11.INIT0 = 16'h5aaa;
    defparam add_215_11.INIT1 = 16'h5aaa;
    defparam add_215_11.INJECT1_0 = "NO";
    defparam add_215_11.INJECT1_1 = "NO";
    FD1S3AY ss_i4_rep_431 (.D(n19947), .CK(clk_N_875), .Q(n22440));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i4_rep_431.GSR = "ENABLED";
    CCU2D add_1188_19 (.A0(n5444), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5446), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18418), 
          .COUT(n18419), .S0(n2353[17]), .S1(n2353[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1188_19.INIT0 = 16'hf555;
    defparam add_1188_19.INIT1 = 16'hf555;
    defparam add_1188_19.INJECT1_0 = "NO";
    defparam add_1188_19.INJECT1_1 = "NO";
    CCU2D add_215_9 (.A0(Out1[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18432), 
          .COUT(n18433), .S0(n1315[7]), .S1(n1315[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_9.INIT0 = 16'h5aaa;
    defparam add_215_9.INIT1 = 16'h5aaa;
    defparam add_215_9.INJECT1_0 = "NO";
    defparam add_215_9.INJECT1_1 = "NO";
    CCU2D add_215_7 (.A0(Out1[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18431), 
          .COUT(n18432), .S0(n1315[5]), .S1(n1315[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_7.INIT0 = 16'h5aaa;
    defparam add_215_7.INIT1 = 16'h5aaa;
    defparam add_215_7.INJECT1_0 = "NO";
    defparam add_215_7.INJECT1_1 = "NO";
    CCU2D add_215_5 (.A0(Out1[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18430), 
          .COUT(n18431), .S0(n1315[3]), .S1(n1315[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_5.INIT0 = 16'h5aaa;
    defparam add_215_5.INIT1 = 16'h5aaa;
    defparam add_215_5.INJECT1_0 = "NO";
    defparam add_215_5.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_21 (.A0(n2353[19]), .B0(n4409), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18666), .COUT(n18667), .S0(n4456), .S1(n4455));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_21.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_21.INIT1 = 16'h5555;
    defparam sub_16_rep_3_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_19 (.A0(n2353[17]), .B0(n4411), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[18]), .B1(n4410), .C1(GND_net), .D1(GND_net), 
          .CIN(n18665), .COUT(n18666), .S0(n4458), .S1(n4457));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_19.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_19.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_19.INJECT1_1 = "NO";
    CCU2D add_215_3 (.A0(Out1[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18429), 
          .COUT(n18430), .S0(n1315[1]), .S1(n1315[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_3.INIT0 = 16'h5aaa;
    defparam add_215_3.INIT1 = 16'h5aaa;
    defparam add_215_3.INJECT1_0 = "NO";
    defparam add_215_3.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_17 (.A0(n2353[15]), .B0(n4413), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[16]), .B1(n4412), .C1(GND_net), .D1(GND_net), 
          .CIN(n18664), .COUT(n18665), .S0(n4460), .S1(n4459));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_17.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_17.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_17.INJECT1_1 = "NO";
    CCU2D add_15369_17 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18784), .S1(n3756));
    defparam add_15369_17.INIT0 = 16'h5555;
    defparam add_15369_17.INIT1 = 16'h0000;
    defparam add_15369_17.INJECT1_0 = "NO";
    defparam add_15369_17.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_15 (.A0(n2353[13]), .B0(n4415), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[14]), .B1(n4414), .C1(GND_net), .D1(GND_net), 
          .CIN(n18663), .COUT(n18664), .S0(n4462), .S1(n4461));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_15.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_15.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_15.INJECT1_1 = "NO";
    CCU2D add_15369_15 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18783), .COUT(n18784));
    defparam add_15369_15.INIT0 = 16'hf555;
    defparam add_15369_15.INIT1 = 16'hf555;
    defparam add_15369_15.INJECT1_0 = "NO";
    defparam add_15369_15.INJECT1_1 = "NO";
    CCU2D add_15369_13 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18782), .COUT(n18783));
    defparam add_15369_13.INIT0 = 16'hf555;
    defparam add_15369_13.INIT1 = 16'hf555;
    defparam add_15369_13.INJECT1_0 = "NO";
    defparam add_15369_13.INJECT1_1 = "NO";
    CCU2D add_215_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[13]), .B1(n18920), .C1(n18921), .D1(Out1[28]), .COUT(n18429), 
          .S1(n1315[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_1.INIT0 = 16'hF000;
    defparam add_215_1.INIT1 = 16'h56aa;
    defparam add_215_1.INJECT1_0 = "NO";
    defparam add_215_1.INJECT1_1 = "NO";
    CCU2D add_223_17 (.A0(Out3[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18452), 
          .S0(n1357[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_17.INIT0 = 16'h5aaa;
    defparam add_223_17.INIT1 = 16'h0000;
    defparam add_223_17.INJECT1_0 = "NO";
    defparam add_223_17.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_13 (.A0(n2353[11]), .B0(n4417), .C0(GND_net), 
          .D0(GND_net), .A1(n2353[12]), .B1(n4416), .C1(GND_net), .D1(GND_net), 
          .CIN(n18662), .COUT(n18663), .S0(n4464), .S1(n4463));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_13.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_13.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_13.INJECT1_1 = "NO";
    CCU2D add_15369_11 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18781), .COUT(n18782));
    defparam add_15369_11.INIT0 = 16'hf555;
    defparam add_15369_11.INIT1 = 16'hf555;
    defparam add_15369_11.INJECT1_0 = "NO";
    defparam add_15369_11.INJECT1_1 = "NO";
    CCU2D add_211_17 (.A0(Out0[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18428), 
          .S0(n1294[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_17.INIT0 = 16'h5aaa;
    defparam add_211_17.INIT1 = 16'h0000;
    defparam add_211_17.INJECT1_0 = "NO";
    defparam add_211_17.INJECT1_1 = "NO";
    CCU2D add_223_15 (.A0(Out3[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18451), 
          .COUT(n18452), .S0(n1357[13]), .S1(n1357[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_15.INIT0 = 16'h5aaa;
    defparam add_223_15.INIT1 = 16'h5aaa;
    defparam add_223_15.INJECT1_0 = "NO";
    defparam add_223_15.INJECT1_1 = "NO";
    CCU2D add_15369_9 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18780), .COUT(n18781));
    defparam add_15369_9.INIT0 = 16'hf555;
    defparam add_15369_9.INIT1 = 16'h0aaa;
    defparam add_15369_9.INJECT1_0 = "NO";
    defparam add_15369_9.INJECT1_1 = "NO";
    FD1S3AX addOut_2102__i1 (.D(n121[1]), .CK(clk_N_875), .Q(addOut[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i1.GSR = "ENABLED";
    PFUMX i17659 (.BLUT(n21736), .ALUT(n21737), .C0(ss[0]), .Z(n4358));
    PFUMX mux_137_i23 (.BLUT(n585[22]), .ALUT(intgOut3[22]), .C0(n21646), 
          .Z(n615[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX i17655 (.BLUT(n21730), .ALUT(n21731), .C0(ss[1]), .Z(n20384));
    PFUMX mux_137_i24 (.BLUT(n585[23]), .ALUT(intgOut3[23]), .C0(n21646), 
          .Z(n615[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i25 (.BLUT(n585[24]), .ALUT(intgOut3[24]), .C0(n21646), 
          .Z(n615[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i26 (.BLUT(n585[25]), .ALUT(intgOut3[25]), .C0(n21646), 
          .Z(n615[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i27 (.BLUT(n585[26]), .ALUT(intgOut3[26]), .C0(n21646), 
          .Z(n615[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i28 (.BLUT(n585[27]), .ALUT(intgOut3[27]), .C0(n21646), 
          .Z(n615[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i29 (.BLUT(n585[28]), .ALUT(intgOut3[28]), .C0(n21646), 
          .Z(n615[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1S3AX addOut_2102__i2 (.D(n121[2]), .CK(clk_N_875), .Q(addOut[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i2.GSR = "ENABLED";
    FD1S3AX addOut_2102__i3 (.D(n121[3]), .CK(clk_N_875), .Q(addOut[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i3.GSR = "ENABLED";
    FD1S3AX addOut_2102__i4 (.D(n121[4]), .CK(clk_N_875), .Q(addOut[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i4.GSR = "ENABLED";
    FD1S3AX addOut_2102__i5 (.D(n121[5]), .CK(clk_N_875), .Q(addOut[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i5.GSR = "ENABLED";
    FD1S3AX addOut_2102__i6 (.D(n121[6]), .CK(clk_N_875), .Q(addOut[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i6.GSR = "ENABLED";
    FD1S3AX addOut_2102__i7 (.D(n121[7]), .CK(clk_N_875), .Q(addOut[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i7.GSR = "ENABLED";
    FD1S3AX addOut_2102__i8 (.D(n121[8]), .CK(clk_N_875), .Q(addOut[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i8.GSR = "ENABLED";
    FD1S3AX addOut_2102__i9 (.D(n121[9]), .CK(clk_N_875), .Q(addOut[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i9.GSR = "ENABLED";
    FD1S3AX addOut_2102__i10 (.D(n121[10]), .CK(clk_N_875), .Q(addOut[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i10.GSR = "ENABLED";
    FD1S3AX addOut_2102__i11 (.D(n121[11]), .CK(clk_N_875), .Q(addOut[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i11.GSR = "ENABLED";
    FD1S3AX addOut_2102__i12 (.D(n121[12]), .CK(clk_N_875), .Q(addOut[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i12.GSR = "ENABLED";
    FD1S3AX addOut_2102__i13 (.D(n121[13]), .CK(clk_N_875), .Q(addOut[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i13.GSR = "ENABLED";
    FD1S3AX addOut_2102__i14 (.D(n121[14]), .CK(clk_N_875), .Q(addOut[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i14.GSR = "ENABLED";
    FD1S3AX addOut_2102__i15 (.D(n121[15]), .CK(clk_N_875), .Q(addOut[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i15.GSR = "ENABLED";
    FD1S3AX addOut_2102__i16 (.D(n121[16]), .CK(clk_N_875), .Q(addOut[16])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i16.GSR = "ENABLED";
    FD1S3AX addOut_2102__i17 (.D(n121[17]), .CK(clk_N_875), .Q(addOut[17])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i17.GSR = "ENABLED";
    FD1S3AX addOut_2102__i18 (.D(n121[18]), .CK(clk_N_875), .Q(addOut[18])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i18.GSR = "ENABLED";
    FD1S3AX addOut_2102__i19 (.D(n121[19]), .CK(clk_N_875), .Q(addOut[19])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i19.GSR = "ENABLED";
    FD1S3AX addOut_2102__i20 (.D(n121[20]), .CK(clk_N_875), .Q(addOut[20])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i20.GSR = "ENABLED";
    FD1S3AX addOut_2102__i21 (.D(n121[21]), .CK(clk_N_875), .Q(addOut[21])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i21.GSR = "ENABLED";
    FD1S3AX addOut_2102__i22 (.D(n121[22]), .CK(clk_N_875), .Q(addOut[22])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i22.GSR = "ENABLED";
    FD1S3AX addOut_2102__i23 (.D(n121[23]), .CK(clk_N_875), .Q(addOut[23])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i23.GSR = "ENABLED";
    FD1S3AX addOut_2102__i24 (.D(n121[24]), .CK(clk_N_875), .Q(addOut[24])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i24.GSR = "ENABLED";
    FD1S3AX addOut_2102__i25 (.D(n121[25]), .CK(clk_N_875), .Q(addOut[25])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i25.GSR = "ENABLED";
    FD1S3AX addOut_2102__i26 (.D(n121[26]), .CK(clk_N_875), .Q(addOut[26])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i26.GSR = "ENABLED";
    FD1S3AX addOut_2102__i27 (.D(n121[27]), .CK(clk_N_875), .Q(addOut[27])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i27.GSR = "ENABLED";
    FD1S3AX addOut_2102__i28 (.D(n121[28]), .CK(clk_N_875), .Q(addOut[28])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2102__i28.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR
//

module PWMGENERATOR (pwm_clk, PWM_m4, free_m4, clkout_c_enable_341, 
            PWMdut_m4, GND_net, hallsense_m4, n21696, enable_m4, n3244, 
            n21700, n3208);
    input pwm_clk;
    output PWM_m4;
    output free_m4;
    input clkout_c_enable_341;
    input [9:0]PWMdut_m4;
    input GND_net;
    input [2:0]hallsense_m4;
    output n21696;
    input enable_m4;
    output n3244;
    output n21700;
    output n3208;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    
    wire n14147;
    wire [9:0]n45;
    
    wire PWM_N_2176, free_N_2188, n17, n16, n10, n7, n10_adj_2325, 
        n11442, n9, n3896, n14, n10_adj_2326, n18512, n18511, 
        n18510, n18509, n18508, n18560, n18559, n18558, n18557, 
        n18556;
    
    FD1S3IX cnt_2106__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14147), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i0.GSR = "ENABLED";
    FD1S3AX PWM_20 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m4)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_2188), .SP(clkout_c_enable_341), .CK(pwm_clk), 
            .Q(free_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i17485_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n14147)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17485_4_lut.init = 16'h0400;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i6_4_lut (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut.init = 16'hffef;
    LUT4 i2_3_lut (.A(PWMdut_m4[5]), .B(PWMdut_m4[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_2325), .B(PWMdut_m4[9]), .C(PWMdut_m4[8]), 
         .D(PWMdut_m4[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2326_3_lut (.A(n11442), .B(PWMdut_m4[4]), .C(PWMdut_m4[3]), 
         .Z(n10_adj_2325)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2326_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1810_1_lut (.A(n3896), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1810_1_lut.init = 16'h5555;
    LUT4 i17463_4_lut (.A(PWMdut_m4[5]), .B(n14), .C(n10_adj_2326), .D(PWMdut_m4[8]), 
         .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17463_4_lut.init = 16'h0001;
    LUT4 i6_4_lut_adj_40 (.A(PWMdut_m4[9]), .B(PWMdut_m4[3]), .C(PWMdut_m4[4]), 
         .D(n11442), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut_adj_40.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[7]), .Z(n10_adj_2326)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_41 (.A(PWMdut_m4[2]), .B(PWMdut_m4[1]), .C(PWMdut_m4[0]), 
         .Z(n11442)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_41.init = 16'hfefe;
    CCU2D sub_1808_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m4[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18512), .S1(n3896));
    defparam sub_1808_add_2_11.INIT0 = 16'h5999;
    defparam sub_1808_add_2_11.INIT1 = 16'h0000;
    defparam sub_1808_add_2_11.INJECT1_0 = "NO";
    defparam sub_1808_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_9 (.A0(PWMdut_m4[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m4[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18511), 
          .COUT(n18512));
    defparam sub_1808_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1808_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1808_add_2_9.INJECT1_0 = "NO";
    defparam sub_1808_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_7 (.A0(PWMdut_m4[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m4[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18510), 
          .COUT(n18511));
    defparam sub_1808_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1808_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1808_add_2_7.INJECT1_0 = "NO";
    defparam sub_1808_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_5 (.A0(PWMdut_m4[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m4[4]), .C1(n9), .D1(n10), .CIN(n18509), 
          .COUT(n18510));
    defparam sub_1808_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1808_add_2_5.INIT1 = 16'h5999;
    defparam sub_1808_add_2_5.INJECT1_0 = "NO";
    defparam sub_1808_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m4[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m4[2]), .C1(n9), .D1(n10), .CIN(n18508), 
          .COUT(n18509));
    defparam sub_1808_add_2_3.INIT0 = 16'h5999;
    defparam sub_1808_add_2_3.INIT1 = 16'h5999;
    defparam sub_1808_add_2_3.INJECT1_0 = "NO";
    defparam sub_1808_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m4[0]), .C1(n9), .D1(n10), 
          .COUT(n18508));
    defparam sub_1808_add_2_1.INIT0 = 16'h0000;
    defparam sub_1808_add_2_1.INIT1 = 16'h5999;
    defparam sub_1808_add_2_1.INJECT1_0 = "NO";
    defparam sub_1808_add_2_1.INJECT1_1 = "NO";
    LUT4 i1722_3_lut_rep_383 (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .Z(n21696)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1722_3_lut_rep_383.init = 16'h1414;
    LUT4 i17535_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .D(enable_m4), .Z(n3244)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17535_2_lut_4_lut.init = 16'hebff;
    LUT4 i1692_3_lut_rep_387 (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .Z(n21700)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1692_3_lut_rep_387.init = 16'h1414;
    LUT4 i17531_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .D(enable_m4), .Z(n3208)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17531_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2106__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14147), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i1.GSR = "ENABLED";
    FD1S3IX cnt_2106__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14147), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i2.GSR = "ENABLED";
    FD1S3IX cnt_2106__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14147), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i3.GSR = "ENABLED";
    FD1S3IX cnt_2106__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14147), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i4.GSR = "ENABLED";
    FD1S3IX cnt_2106__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14147), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i5.GSR = "ENABLED";
    FD1S3IX cnt_2106__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14147), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i6.GSR = "ENABLED";
    FD1S3IX cnt_2106__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14147), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i7.GSR = "ENABLED";
    FD1S3IX cnt_2106__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14147), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i8.GSR = "ENABLED";
    FD1S3IX cnt_2106__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14147), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106__i9.GSR = "ENABLED";
    CCU2D cnt_2106_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18560), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2106_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2106_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2106_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2106_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18559), 
          .COUT(n18560), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2106_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2106_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2106_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2106_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18558), 
          .COUT(n18559), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2106_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2106_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2106_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2106_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18557), 
          .COUT(n18558), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2106_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2106_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2106_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2106_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18556), 
          .COUT(n18557), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2106_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2106_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2106_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2106_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18556), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2106_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2106_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2106_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2106_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module HALL
//

module HALL (clk_1mhz, \speed_m4[0] , hallsense_m4, clkout_c_enable_272, 
            clkout_c_enable_341, H_A_m4_c, H_B_m4_c, H_C_m4_c, \speed_m4[1] , 
            \speed_m4[2] , \speed_m4[3] , \speed_m4[4] , \speed_m4[5] , 
            \speed_m4[6] , \speed_m4[7] , \speed_m4[8] , \speed_m4[9] , 
            \speed_m4[10] , \speed_m4[11] , \speed_m4[12] , \speed_m4[13] , 
            \speed_m4[14] , \speed_m4[15] , \speed_m4[16] , \speed_m4[17] , 
            \speed_m4[18] , \speed_m4[19] , GND_net, n22430);
    input clk_1mhz;
    output \speed_m4[0] ;
    output [2:0]hallsense_m4;
    input clkout_c_enable_272;
    input clkout_c_enable_341;
    input H_A_m4_c;
    input H_B_m4_c;
    input H_C_m4_c;
    output \speed_m4[1] ;
    output \speed_m4[2] ;
    output \speed_m4[3] ;
    output \speed_m4[4] ;
    output \speed_m4[5] ;
    output \speed_m4[6] ;
    output \speed_m4[7] ;
    output \speed_m4[8] ;
    output \speed_m4[9] ;
    output \speed_m4[10] ;
    output \speed_m4[11] ;
    output \speed_m4[12] ;
    output \speed_m4[13] ;
    output \speed_m4[14] ;
    output \speed_m4[15] ;
    output \speed_m4[16] ;
    output \speed_m4[17] ;
    output \speed_m4[18] ;
    output \speed_m4[19] ;
    input GND_net;
    input n22430;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21720;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_89;
    wire [19:0]count_19__N_2067;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4605, stable_counting;
    wire [19:0]speedt_19__N_2047;
    
    wire hall3_lat, hall3_old, hall1_lat, n21679, n21643, n4, n19077, 
        n20024, clk_1mhz_enable_185, hall2_lat, n21, n19839, n26, 
        n22, hall1_old, hall2_old, n19992, n21718, n21719, n19986;
    wire [6:0]n63;
    
    wire n11458, n11451, stable_counting_N_2129, n20190, n21717, n20172, 
        n20060, n20124, n19934, n21653, n19811, n21639, n4_adj_2324, 
        n21652, n21680, n14393, n18492, n18491, n18490, n21663, 
        n18489, n18488, n18487, n18486, n18485, n18484, n18483;
    
    LUT4 i2539_2_lut_rep_407 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21720)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2539_2_lut_rep_407.init = 16'h8888;
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2067[0]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_19__N_2067[0]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_2047[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_272), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m4_c), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    LUT4 i2565_2_lut_rep_330_3_lut_4_lut (.A(stable_count[3]), .B(n21679), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21643)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2565_2_lut_rep_330_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21679), .C(stable_count[0]), 
         .D(stable_count[4]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i17558_4_lut (.A(n19077), .B(n20024), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_185)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17558_4_lut.init = 16'hdffd;
    FD1P3AX hall2_lat_58 (.D(H_B_m4_c), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n21), .B(n19839), .C(n26), .D(n22), .Z(n19077)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i16627_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n20024)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16627_4_lut.init = 16'h7bde;
    LUT4 i12_4_lut (.A(n19992), .B(n21718), .C(n21719), .D(n19986), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[11]), .B(count[7]), .C(count[16]), .D(count[17]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i8_4_lut.init = 16'hfffe;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    LUT4 i2535_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2535_1_lut.init = 16'h5555;
    FD1P3AX hall3_lat_59 (.D(H_C_m4_c), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_341), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 i11516_4_lut (.A(n11458), .B(n11451), .C(stable_counting), .D(stable_counting_N_2129), 
         .Z(clk_1mhz_enable_89)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11516_4_lut.init = 16'hcaea;
    LUT4 i4_4_lut (.A(count[8]), .B(n20190), .C(n19839), .D(n21717), 
         .Z(n11458)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h2000;
    LUT4 i16792_4_lut (.A(n19986), .B(n20172), .C(count[6]), .D(n20060), 
         .Z(n20190)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16792_4_lut.init = 16'hfffe;
    LUT4 i16774_4_lut (.A(count[11]), .B(n20124), .C(n19992), .D(count[7]), 
         .Z(n20172)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16774_4_lut.init = 16'hfffe;
    LUT4 i16663_2_lut (.A(count[16]), .B(count[17]), .Z(n20060)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16663_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(n19934), .B(stable_count[0]), .C(n21653), .D(n19811), 
         .Z(n11451)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_adj_37 (.A(n63[2]), .B(n19934), .C(n21639), .D(n4), 
         .Z(stable_counting_N_2129)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_37.init = 16'h0004;
    LUT4 i1_4_lut_adj_38 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4_adj_2324)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_38.init = 16'h7bde;
    LUT4 i2537_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2537_2_lut.init = 16'h6666;
    LUT4 i16595_2_lut (.A(count[4]), .B(count[5]), .Z(n19992)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16595_2_lut.init = 16'heeee;
    LUT4 i16589_2_lut (.A(count[18]), .B(count[15]), .Z(n19986)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16589_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(count[9]), .B(count[0]), .C(count[2]), .D(count[10]), 
         .Z(n19839)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2047[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2047[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2047[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2047[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2047[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2047[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2047[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2047[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2047[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2047[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2047[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2047[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2067[1]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2067[2]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2067[3]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2067[4]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2067[5]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2067[6]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2067[7]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2067[8]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2067[9]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2067[10]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2067[11]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2067[12]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2067[13]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2067[14]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2067[15]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2067[16]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2067[17]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2067[18]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2067[19]), .SP(clk_1mhz_enable_89), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2047[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2047[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2047[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX count__i1 (.D(count_19__N_2067[1]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2067[2]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2067[3]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2067[4]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2067[5]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2067[6]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2067[7]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2067[8]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2067[9]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2067[10]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2067[11]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2067[12]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2067[13]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2067[14]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2067[15]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2067[16]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2067[17]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2067[18]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2067[19]), .CK(clk_1mhz), .CD(n4605), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3AX speed__i2 (.D(speedt_19__N_2047[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2047[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2047[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2047[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2047[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2047[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2047[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2047[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2047[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2047[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2047[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2047[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2047[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2047[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2047[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2047[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2047[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2047[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2047[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2047[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2047[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2047[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2047[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11458), .B(n11451), .C(count_19__N_2067[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2047[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2278_2_lut (.A(stable_counting), .B(stable_counting_N_2129), .Z(n4605)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2278_2_lut.init = 16'h8888;
    LUT4 i2560_2_lut_rep_339_3_lut_4_lut (.A(stable_count[2]), .B(n21720), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21652)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2560_2_lut_rep_339_3_lut_4_lut.init = 16'h8000;
    LUT4 i2558_2_lut_rep_340_3_lut_4_lut (.A(stable_count[2]), .B(n21720), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21653)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2558_2_lut_rep_340_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2_3_lut_rep_367 (.A(hall3_old), .B(n4_adj_2324), .C(hall3_lat), 
         .Z(n21680)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_367.init = 16'hdede;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4_adj_2324), .C(hall3_lat), 
         .D(n63[1]), .Z(n19934)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 i1_2_lut_4_lut_adj_39 (.A(n63[3]), .B(n63[6]), .C(n21643), .D(n63[2]), 
         .Z(n19811)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_39.init = 16'hfffe;
    LUT4 i2_3_lut_rep_326_4_lut (.A(stable_count[5]), .B(n21652), .C(n63[6]), 
         .D(n63[3]), .Z(n21639)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_326_4_lut.init = 16'hfff6;
    LUT4 i2544_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2544_2_lut_3_lut.init = 16'h7878;
    LUT4 i16746_3_lut (.A(n21680), .B(stable_counting), .C(stable_counting_N_2129), 
         .Z(n14393)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16746_3_lut.init = 16'hc8c8;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21643), .SP(stable_counting), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21653), .SP(stable_counting), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18492), 
          .S0(count_19__N_2067[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18491), .COUT(n18492), .S0(count_19__N_2067[17]), .S1(count_19__N_2067[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18490), .COUT(n18491), .S0(count_19__N_2067[15]), .S1(count_19__N_2067[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    FD1P3IX stable_counting_62 (.D(n22430), .SP(clk_1mhz_enable_185), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14393), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    LUT4 i16704_2_lut_rep_404 (.A(count[3]), .B(count[13]), .Z(n21717)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16704_2_lut_rep_404.init = 16'h8888;
    LUT4 i16593_2_lut_rep_406 (.A(count[12]), .B(count[19]), .Z(n21719)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16593_2_lut_rep_406.init = 16'heeee;
    LUT4 i16726_2_lut_3_lut_4_lut (.A(count[12]), .B(count[19]), .C(count[1]), 
         .D(count[14]), .Z(n20124)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16726_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2551_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2551_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i16591_2_lut_rep_405 (.A(count[14]), .B(count[1]), .Z(n21718)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16591_2_lut_rep_405.init = 16'heeee;
    LUT4 i2546_2_lut_rep_366_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21679)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2546_2_lut_rep_366_3_lut.init = 16'h8080;
    LUT4 i2553_2_lut_rep_350_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21663)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2553_2_lut_rep_350_3_lut_4_lut.init = 16'h8000;
    LUT4 i7_3_lut_4_lut (.A(count[3]), .B(count[13]), .C(count[8]), .D(count[6]), 
         .Z(n21)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i7_3_lut_4_lut.init = 16'hff7f;
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18489), .COUT(n18490), .S0(count_19__N_2067[13]), .S1(count_19__N_2067[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    LUT4 i2572_3_lut_4_lut (.A(stable_count[4]), .B(n21663), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2572_3_lut_4_lut.init = 16'h7f80;
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18488), .COUT(n18489), .S0(count_19__N_2067[11]), .S1(count_19__N_2067[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18487), .COUT(n18488), .S0(count_19__N_2067[9]), .S1(count_19__N_2067[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18486), 
          .COUT(n18487), .S0(count_19__N_2067[7]), .S1(count_19__N_2067[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18485), 
          .COUT(n18486), .S0(count_19__N_2067[5]), .S1(count_19__N_2067[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18484), 
          .COUT(n18485), .S0(count_19__N_2067[3]), .S1(count_19__N_2067[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18483), 
          .COUT(n18484), .S0(count_19__N_2067[1]), .S1(count_19__N_2067[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18483), 
          .S1(count_19__N_2067[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    
endmodule
