// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.8.0.115.3
// Netlist written on Mon May 22 15:05:12 2017
//
// Verilog Description of module SPI_loopback_Top
//

module SPI_loopback_Top (CS, SCK, MOSI, MISO, HALL_A_OUT, HALL_B_OUT, 
            HALL_C_OUT, LED1, LED2, LED3, LED4, clkout, H_A_m1, 
            H_B_m1, H_C_m1, MA_m1, MB_m1, MC_m1, H_A_m2, H_B_m2, 
            H_C_m2, MA_m2, MB_m2, MC_m2, H_A_m3, H_B_m3, H_C_m3, 
            MA_m3, MB_m3, MC_m3, H_A_m4, H_B_m4, H_C_m4, MA_m4, 
            MB_m4, MC_m4);   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(24[8:24])
    input CS;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(27[2:4])
    input SCK;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(28[2:5])
    input MOSI;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(29[2:6])
    output MISO;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(30[2:6])
    output HALL_A_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(33[2:12])
    output HALL_B_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(34[2:12])
    output HALL_C_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(35[2:12])
    output LED1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(38[2:6])
    output LED2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(39[2:6])
    output LED3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(40[2:6])
    output LED4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(41[2:6])
    output clkout;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    input H_A_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(47[2:8])
    input H_B_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(48[2:8])
    input H_C_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(49[2:8])
    output [1:0]MA_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    output [1:0]MB_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    output [1:0]MC_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    input H_A_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(55[2:8])
    input H_B_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(56[2:8])
    input H_C_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(57[2:8])
    output [1:0]MA_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    output [1:0]MB_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    output [1:0]MC_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    input H_A_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(63[2:8])
    input H_B_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(64[2:8])
    input H_C_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(65[2:8])
    output [1:0]MA_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    output [1:0]MB_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    output [1:0]MC_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    input H_A_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(71[2:8])
    input H_B_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(72[2:8])
    input H_C_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(73[2:8])
    output [1:0]MA_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    output [1:0]MB_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    output [1:0]MC_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    
    wire GND_net, VCC_net, CS_c, SCK_c, MOSI_c, HALL_A_OUT_c_c, 
        HALL_B_OUT_c_c, HALL_C_OUT_c_c, LED1_c, LED2_c, LED3_c, LED4_c, 
        H_A_m1_c, H_B_m1_c, H_C_m1_c, MA_m1_c_1, MA_m1_c_0, MB_m1_c_1, 
        MB_m1_c_0, MC_m1_c_1, MC_m1_c_0, H_A_m2_c, H_B_m2_c, H_C_m2_c, 
        MA_m2_c_1, MA_m2_c_0, MB_m2_c_1, MB_m2_c_0, MC_m2_c_1, MC_m2_c_0, 
        H_A_m3_c, H_B_m3_c, H_C_m3_c, MA_m3_c_1, MA_m3_c_0, MB_m3_c_1, 
        MB_m3_c_0, MC_m3_c_1, MC_m3_c_0, MA_m4_c_1, MA_m4_c_0, MB_m4_c_1, 
        MB_m4_c_0, MC_m4_c_1, MC_m4_c_0, rst, enable_m1, enable_m2, 
        enable_m3, enable_m4;
    wire [20:0]speed_set_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(99[9:21])
    wire [20:0]speed_set_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(100[9:21])
    wire [20:0]speed_set_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(101[9:21])
    wire [20:0]speed_set_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(102[9:21])
    wire [20:0]speed_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(104[9:17])
    wire [20:0]speed_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(105[9:17])
    wire [20:0]speed_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(106[9:17])
    wire [20:0]speed_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(107[9:17])
    wire [2:0]hallsense_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(110[9:21])
    wire [2:0]hallsense_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(111[9:21])
    wire [2:0]hallsense_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(112[9:21])
    wire [2:0]hallsense_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(113[9:21])
    
    wire PWM_m1, PWM_m2, PWM_m3, PWM_m4;
    wire [9:0]PWMdut_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(120[9:18])
    wire [9:0]PWMdut_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(121[9:18])
    wire [9:0]PWMdut_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(122[9:18])
    wire [9:0]PWMdut_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(123[9:18])
    
    wire dir_m1, dir_m2, dir_m3, dir_m4;
    wire [13:0]start_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(135[9:18])
    
    wire free_m1, free_m2, free_m3, free_m4;
    wire [20:0]speed_avg_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(144[9:21])
    wire [20:0]speed_avg_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(145[9:21])
    wire [20:0]speed_avg_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(146[9:21])
    wire [20:0]speed_avg_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(147[9:21])
    wire [95:0]send_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(67[10:21])
    
    wire n22100, n75, n74, n73, n72, n71, n70, n69, n68, n67, 
        n66, n65, n64, n63, n62, n3278, n3220, n3184, n3232, 
        n3196, n3170, n3112, n3076, n3124, n3088, n3062, n3004;
    wire [95:0]send_buffer_95__N_346;
    
    wire n2968, n3016, n2980, n2954, n2896, MISO_N_624, n4434, 
        n18445, n2872;
    wire [25:0]subOut_24__N_1177;
    
    wire n19411, n2860, n4461, n4458, n4455, n4452, n4435, n4447, 
        n4430, n4427, n4425, n4422, n4417, n4414, n5, n7, n3, 
        n18510, n20284, n19427, n18938, n19415, n21328, n22097, 
        n2908, n4322, n4448, n4446, n4445, n4444, n4443, n4442, 
        n4441, n4440, n4436, n4433, n4432, n4431, n4429, n4428, 
        n4426, n4424, n4423, n4421, n4420, n4419, n4418, n4416, 
        n4415, n18509, n4460, n4459, n4457, n4456, n4454, n4453, 
        n4451, n4450, n4449, n5132, n10392, n6, n19421, n21309, 
        n18181, n18180, n18179, n18178, n18177, n18176, n18175, 
        clkout_c_enable_173, clkout_c_enable_266, clkout_c_enable_172, 
        n21375, n21373, n21372, n21371, n21369, n21368, n21366, 
        n21363, n21362, n21361, n21358, n21357, n21354, n21336;
    
    VHI i2 (.Z(VCC_net));
    OSCH OSCInst0 (.STDBY(GND_net), .OSC(clkout_c)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCInst0.NOM_FREQ = "38.00";
    LUT4 i13066_4_lut (.A(n4322), .B(speed_avg_m3[19]), .C(n21328), .D(speed_avg_m4[19]), 
         .Z(n3)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i13066_4_lut.init = 16'hcac0;
    LUT4 mux_2142_i1_3_lut (.A(n4436), .B(n4461), .C(n18938), .Z(subOut_24__N_1177[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i1_3_lut.init = 16'hacac;
    LUT4 m1_lut (.Z(n22097)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    OB MA_m2_pad_0 (.I(MA_m2_c_0), .O(MA_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    LUT4 i1_2_lut_4_lut (.A(send_buffer[94]), .B(speed_avg_m1[19]), .C(n21354), 
         .D(n21336), .Z(send_buffer_95__N_346[94])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(73[10:15])
    defparam i1_2_lut_4_lut.init = 16'h00ca;
    FD1P3AX start_cnt_2076__i0 (.D(n75), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i0.GSR = "DISABLED";
    LUT4 mux_2142_i21_3_lut (.A(n4416), .B(n4441), .C(n18938), .Z(subOut_24__N_1177[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i21_3_lut.init = 16'hacac;
    OB HALL_B_OUT_pad (.I(HALL_B_OUT_c_c), .O(HALL_B_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(34[2:12])
    OB HALL_A_OUT_pad (.I(HALL_A_OUT_c_c), .O(HALL_A_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(33[2:12])
    OB MA_m2_pad_1 (.I(MA_m2_c_1), .O(MA_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    IB H_B_m1_pad (.I(H_B_m1), .O(H_B_m1_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(48[2:8])
    OBZ n5131_pad (.I(MISO_N_624), .T(n5132), .O(MISO));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    IB H_A_m1_pad (.I(H_A_m1), .O(H_A_m1_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(47[2:8])
    IB MOSI_pad (.I(MOSI), .O(MOSI_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(29[2:6])
    IB SCK_pad (.I(SCK), .O(SCK_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(28[2:5])
    IB CS_pad (.I(CS), .O(CS_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(27[2:4])
    OB MC_m4_pad_0 (.I(MC_m4_c_0), .O(MC_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    OB MC_m4_pad_1 (.I(MC_m4_c_1), .O(MC_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    OB MB_m4_pad_0 (.I(MB_m4_c_0), .O(MB_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    OB MB_m4_pad_1 (.I(MB_m4_c_1), .O(MB_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    OB MC_m1_pad_0 (.I(MC_m1_c_0), .O(MC_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    OB MC_m1_pad_1 (.I(MC_m1_c_1), .O(MC_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    OB MA_m4_pad_0 (.I(MA_m4_c_0), .O(MA_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_0 (.I(MB_m1_c_0), .O(MB_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    OB MA_m4_pad_1 (.I(MA_m4_c_1), .O(MA_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_1 (.I(MB_m1_c_1), .O(MB_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    OB MC_m3_pad_0 (.I(MC_m3_c_0), .O(MC_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    IB HALL_C_OUT_c_pad (.I(H_C_m4), .O(HALL_C_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(73[2:8])
    OB MA_m1_pad_0 (.I(MA_m1_c_0), .O(MA_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    OB MC_m3_pad_1 (.I(MC_m3_c_1), .O(MC_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    IB HALL_B_OUT_c_pad (.I(H_B_m4), .O(HALL_B_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(72[2:8])
    OB MA_m1_pad_1 (.I(MA_m1_c_1), .O(MA_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    OB MB_m3_pad_0 (.I(MB_m3_c_0), .O(MB_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    IB HALL_A_OUT_c_pad (.I(H_A_m4), .O(HALL_A_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(71[2:8])
    OB clkout_pad (.I(clkout_c), .O(clkout));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    OB MB_m3_pad_1 (.I(MB_m3_c_1), .O(MB_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    IB H_C_m3_pad (.I(H_C_m3), .O(H_C_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(65[2:8])
    OB LED4_pad (.I(LED4_c), .O(LED4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(41[2:6])
    OB MA_m3_pad_0 (.I(MA_m3_c_0), .O(MA_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    IB H_B_m3_pad (.I(H_B_m3), .O(H_B_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(64[2:8])
    OB LED3_pad (.I(LED3_c), .O(LED3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(40[2:6])
    OB MA_m3_pad_1 (.I(MA_m3_c_1), .O(MA_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    IB H_A_m3_pad (.I(H_A_m3), .O(H_A_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(63[2:8])
    OB LED2_pad (.I(LED2_c), .O(LED2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(39[2:6])
    OB MC_m2_pad_0 (.I(MC_m2_c_0), .O(MC_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    IB H_C_m2_pad (.I(H_C_m2), .O(H_C_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(57[2:8])
    OB LED1_pad (.I(LED1_c), .O(LED1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(38[2:6])
    OB MC_m2_pad_1 (.I(MC_m2_c_1), .O(MC_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    IB H_B_m2_pad (.I(H_B_m2), .O(H_B_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(56[2:8])
    OB HALL_C_OUT_pad (.I(HALL_C_OUT_c_c), .O(HALL_C_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(35[2:12])
    OB MB_m2_pad_0 (.I(MB_m2_c_0), .O(MB_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    IB H_A_m2_pad (.I(H_A_m2), .O(H_A_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(55[2:8])
    OB MB_m2_pad_1 (.I(MB_m2_c_1), .O(MB_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    IB H_C_m1_pad (.I(H_C_m1), .O(H_C_m1_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(49[2:8])
    FD1S3AX rst_12_rep_411 (.D(n21309), .CK(clkout_c), .Q(clkout_c_enable_173));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12_rep_411.GSR = "DISABLED";
    FD1S3AX rst_12_rep_410 (.D(n21309), .CK(clkout_c), .Q(clkout_c_enable_172));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12_rep_410.GSR = "DISABLED";
    CCU2D start_cnt_2076_add_4_15 (.A0(start_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18181), .S0(n62));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_15.INIT0 = 16'hfaaa;
    defparam start_cnt_2076_add_4_15.INIT1 = 16'h0000;
    defparam start_cnt_2076_add_4_15.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_15.INJECT1_1 = "NO";
    CCU2D start_cnt_2076_add_4_13 (.A0(start_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18180), .COUT(n18181), .S0(n64), .S1(n63));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_13.INIT0 = 16'hfaaa;
    defparam start_cnt_2076_add_4_13.INIT1 = 16'hfaaa;
    defparam start_cnt_2076_add_4_13.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_13.INJECT1_1 = "NO";
    CCU2D start_cnt_2076_add_4_11 (.A0(start_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18179), .COUT(n18180), .S0(n66), .S1(n65));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_11.INIT0 = 16'hfaaa;
    defparam start_cnt_2076_add_4_11.INIT1 = 16'hfaaa;
    defparam start_cnt_2076_add_4_11.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_11.INJECT1_1 = "NO";
    CCU2D start_cnt_2076_add_4_9 (.A0(start_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18178), .COUT(n18179), .S0(n68), .S1(n67));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_9.INIT0 = 16'hfaaa;
    defparam start_cnt_2076_add_4_9.INIT1 = 16'hfaaa;
    defparam start_cnt_2076_add_4_9.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_9.INJECT1_1 = "NO";
    CCU2D start_cnt_2076_add_4_7 (.A0(start_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18177), .COUT(n18178), .S0(n70), .S1(n69));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_7.INIT0 = 16'hfaaa;
    defparam start_cnt_2076_add_4_7.INIT1 = 16'hfaaa;
    defparam start_cnt_2076_add_4_7.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_7.INJECT1_1 = "NO";
    CCU2D start_cnt_2076_add_4_5 (.A0(start_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18176), .COUT(n18177), .S0(n72), .S1(n71));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_5.INIT0 = 16'hfaaa;
    defparam start_cnt_2076_add_4_5.INIT1 = 16'hfaaa;
    defparam start_cnt_2076_add_4_5.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_5.INJECT1_1 = "NO";
    CCU2D start_cnt_2076_add_4_3 (.A0(start_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18175), .COUT(n18176), .S0(n74), .S1(n73));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_3.INIT0 = 16'hfaaa;
    defparam start_cnt_2076_add_4_3.INIT1 = 16'hfaaa;
    defparam start_cnt_2076_add_4_3.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_3.INJECT1_1 = "NO";
    CCU2D start_cnt_2076_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18175), .S1(n75));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076_add_4_1.INIT0 = 16'hF000;
    defparam start_cnt_2076_add_4_1.INIT1 = 16'h0555;
    defparam start_cnt_2076_add_4_1.INJECT1_0 = "NO";
    defparam start_cnt_2076_add_4_1.INJECT1_1 = "NO";
    FD1S3AX rst_12 (.D(n21309), .CK(clkout_c), .Q(rst));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12.GSR = "DISABLED";
    GSR GSR_INST (.GSR(n22100));
    LUT4 i3_4_lut (.A(n18510), .B(start_cnt[10]), .C(start_cnt[9]), .D(start_cnt[8]), 
         .Z(n18445)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_177 (.A(n18509), .B(n6), .C(start_cnt[6]), .D(start_cnt[4]), 
         .Z(n18510)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_177.init = 16'hfefc;
    LUT4 i3_4_lut_adj_178 (.A(start_cnt[0]), .B(start_cnt[3]), .C(start_cnt[2]), 
         .D(start_cnt[1]), .Z(n18509)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_178.init = 16'hfffe;
    LUT4 i2_2_lut (.A(start_cnt[7]), .B(start_cnt[5]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1734_3_lut_rep_376 (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .Z(n21357)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i1734_3_lut_rep_376.init = 16'h4242;
    LUT4 i17207_2_lut_4_lut (.A(hallsense_m4[2]), .B(dir_m4), .C(hallsense_m4[0]), 
         .D(free_m4), .Z(n3278)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i17207_2_lut_4_lut.init = 16'hffbd;
    LUT4 mux_2142_i2_3_lut (.A(n4435), .B(n4460), .C(n18938), .Z(subOut_24__N_1177[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i2_3_lut.init = 16'hacac;
    LUT4 mux_2142_i3_3_lut (.A(n4434), .B(n4459), .C(n18938), .Z(subOut_24__N_1177[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i3_3_lut.init = 16'hacac;
    LUT4 i1644_3_lut_rep_381 (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .Z(n21362)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i1644_3_lut_rep_381.init = 16'h4242;
    LUT4 mux_2142_i4_3_lut (.A(n4433), .B(n4458), .C(n18938), .Z(subOut_24__N_1177[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i4_3_lut.init = 16'hacac;
    LUT4 i17209_2_lut_4_lut (.A(hallsense_m3[2]), .B(dir_m3), .C(hallsense_m3[0]), 
         .D(free_m3), .Z(n3170)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i17209_2_lut_4_lut.init = 16'hffbd;
    LUT4 mux_2142_i5_3_lut (.A(n4432), .B(n4457), .C(n18938), .Z(subOut_24__N_1177[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i5_3_lut.init = 16'hacac;
    PFUMX i13070 (.BLUT(n3), .ALUT(n5), .C0(n20284), .Z(n7));
    LUT4 mux_2142_i6_3_lut (.A(n4431), .B(n4456), .C(n18938), .Z(subOut_24__N_1177[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i6_3_lut.init = 16'hacac;
    LUT4 mux_2142_i7_3_lut (.A(n4430), .B(n4455), .C(n18938), .Z(subOut_24__N_1177[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i7_3_lut.init = 16'hacac;
    LUT4 i1554_3_lut_rep_387 (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .Z(n21368)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i1554_3_lut_rep_387.init = 16'h4242;
    LUT4 i17211_2_lut_4_lut (.A(hallsense_m2[2]), .B(dir_m2), .C(hallsense_m2[0]), 
         .D(free_m2), .Z(n3062)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i17211_2_lut_4_lut.init = 16'hffbd;
    LUT4 mux_2142_i8_3_lut (.A(n4429), .B(n4454), .C(n18938), .Z(subOut_24__N_1177[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i8_3_lut.init = 16'hacac;
    COMMUTATION_U6 COM_I_M3 (.MB_m3_c_0(MB_m3_c_0), .clkout_c(clkout_c), 
            .MC_m3_c_0(MC_m3_c_0), .MA_m3_c_0(MA_m3_c_0), .LED3_c(LED3_c), 
            .enable_m3(enable_m3), .n3076(n3076), .n21366(n21366), .PWM_m3(PWM_m3), 
            .n3112(n3112), .n21363(n21363), .n19427(n19427), .n21362(n21362), 
            .free_m3(free_m3), .MA_m3_c_1(MA_m3_c_1), .n3170(n3170), .MC_m3_c_1(MC_m3_c_1), 
            .n3124(n3124), .MB_m3_c_1(MB_m3_c_1), .n3088(n3088));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(339[13:24])
    LUT4 i1464_3_lut_rep_391 (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .Z(n21372)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i1464_3_lut_rep_391.init = 16'h4242;
    LUT4 i17213_2_lut_4_lut (.A(hallsense_m1[2]), .B(dir_m1), .C(hallsense_m1[0]), 
         .D(free_m1), .Z(n2954)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i17213_2_lut_4_lut.init = 16'hffbd;
    COMMUTATION_U7 COM_I_M2 (.MB_m2_c_0(MB_m2_c_0), .clkout_c(clkout_c), 
            .MC_m2_c_0(MC_m2_c_0), .MA_m2_c_0(MA_m2_c_0), .LED2_c(LED2_c), 
            .enable_m2(enable_m2), .n2968(n2968), .n21371(n21371), .PWM_m2(PWM_m2), 
            .n3004(n3004), .n21369(n21369), .n19411(n19411), .n21368(n21368), 
            .free_m2(free_m2), .MA_m2_c_1(MA_m2_c_1), .n3062(n3062), .MC_m2_c_1(MC_m2_c_1), 
            .n3016(n3016), .MB_m2_c_1(MB_m2_c_1), .n2980(n2980));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(329[13:24])
    COMMUTATION_U8 COM_I_M1 (.MB_m1_c_0(MB_m1_c_0), .clkout_c(clkout_c), 
            .MC_m1_c_0(MC_m1_c_0), .MA_m1_c_0(MA_m1_c_0), .LED1_c(LED1_c), 
            .enable_m1(enable_m1), .n2860(n2860), .n21375(n21375), .PWM_m1(PWM_m1), 
            .n2896(n2896), .n21373(n21373), .n19421(n19421), .n21372(n21372), 
            .free_m1(free_m1), .MA_m1_c_1(MA_m1_c_1), .n2954(n2954), .MC_m1_c_1(MC_m1_c_1), 
            .n2908(n2908), .MB_m1_c_1(MB_m1_c_1), .n2872(n2872));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(319[13:24])
    CLKDIV CLKDIV_I (.clkout_c(clkout_c), .clk_1mhz(clk_1mhz), .pwm_clk(pwm_clk), 
           .GND_net(GND_net), .clk_N_683(clk_N_683));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(302[14:20])
    LUT4 mux_2142_i9_3_lut (.A(n4428), .B(n4453), .C(n18938), .Z(subOut_24__N_1177[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i9_3_lut.init = 16'hacac;
    LUT4 mux_2142_i10_3_lut (.A(n4427), .B(n4452), .C(n18938), .Z(subOut_24__N_1177[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i10_3_lut.init = 16'hacac;
    LUT4 mux_2142_i11_3_lut (.A(n4426), .B(n4451), .C(n18938), .Z(subOut_24__N_1177[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i11_3_lut.init = 16'hacac;
    LUT4 mux_2142_i12_3_lut (.A(n4425), .B(n4450), .C(n18938), .Z(subOut_24__N_1177[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i12_3_lut.init = 16'hacac;
    LUT4 mux_2142_i13_3_lut (.A(n4424), .B(n4449), .C(n18938), .Z(subOut_24__N_1177[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i13_3_lut.init = 16'hacac;
    LUT4 mux_2142_i14_3_lut (.A(n4423), .B(n4448), .C(n18938), .Z(subOut_24__N_1177[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i14_3_lut.init = 16'hacac;
    LUT4 mux_2142_i15_3_lut (.A(n4422), .B(n4447), .C(n18938), .Z(subOut_24__N_1177[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i15_3_lut.init = 16'hacac;
    LUT4 mux_2142_i16_3_lut (.A(n4421), .B(n4446), .C(n18938), .Z(subOut_24__N_1177[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i16_3_lut.init = 16'hacac;
    LUT4 mux_2142_i17_3_lut (.A(n4420), .B(n4445), .C(n18938), .Z(subOut_24__N_1177[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i17_3_lut.init = 16'hacac;
    LUT4 mux_2142_i18_3_lut (.A(n4419), .B(n4444), .C(n18938), .Z(subOut_24__N_1177[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i18_3_lut.init = 16'hacac;
    LUT4 mux_2142_i19_3_lut (.A(n4418), .B(n4443), .C(n18938), .Z(subOut_24__N_1177[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i19_3_lut.init = 16'hacac;
    LUT4 mux_2142_i22_3_lut (.A(n4415), .B(n4440), .C(n18938), .Z(subOut_24__N_1177[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i22_3_lut.init = 16'hacac;
    LUT4 mux_2142_i20_3_lut (.A(n4417), .B(n4442), .C(n18938), .Z(subOut_24__N_1177[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i20_3_lut.init = 16'hacac;
    LUT4 mux_2142_i25_3_lut (.A(n4414), .B(n4440), .C(n18938), .Z(subOut_24__N_1177[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2142_i25_3_lut.init = 16'hacac;
    LUT4 i7910_2_lut (.A(n21309), .B(n62), .Z(n10392)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam i7910_2_lut.init = 16'heeee;
    LUT4 i2341_4_lut_rep_328 (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18445), .Z(n21309)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2341_4_lut_rep_328.init = 16'hccc8;
    LUT4 i9295_1_lut_4_lut (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18445), .Z(clkout_c_enable_266)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i9295_1_lut_4_lut.init = 16'h3337;
    COMMUTATION COM_I_M4 (.MB_m4_c_0(MB_m4_c_0), .clkout_c(clkout_c), .MC_m4_c_0(MC_m4_c_0), 
            .MA_m4_c_0(MA_m4_c_0), .LED4_c(LED4_c), .enable_m4(enable_m4), 
            .n3184(n3184), .n21361(n21361), .PWM_m4(PWM_m4), .n3220(n3220), 
            .n21358(n21358), .n19415(n19415), .n21357(n21357), .free_m4(free_m4), 
            .MA_m4_c_1(MA_m4_c_1), .n3278(n3278), .MC_m4_c_1(MC_m4_c_1), 
            .n3232(n3232), .MB_m4_c_1(MB_m4_c_1), .n3196(n3196));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(349[13:24])
    HALL_U4 HALL_I_M2 (.clk_1mhz(clk_1mhz), .n22097(n22097), .\speed_m2[0] (speed_m2[0]), 
            .hallsense_m2({hallsense_m2}), .clkout_c_enable_173(clkout_c_enable_173), 
            .H_C_m2_c(H_C_m2_c), .rst(rst), .H_A_m2_c(H_A_m2_c), .H_B_m2_c(H_B_m2_c), 
            .\speed_m2[1] (speed_m2[1]), .\speed_m2[2] (speed_m2[2]), .\speed_m2[3] (speed_m2[3]), 
            .\speed_m2[4] (speed_m2[4]), .\speed_m2[5] (speed_m2[5]), .\speed_m2[6] (speed_m2[6]), 
            .\speed_m2[7] (speed_m2[7]), .\speed_m2[8] (speed_m2[8]), .\speed_m2[9] (speed_m2[9]), 
            .\speed_m2[10] (speed_m2[10]), .\speed_m2[11] (speed_m2[11]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_m2[13] (speed_m2[13]), 
            .\speed_m2[14] (speed_m2[14]), .\speed_m2[15] (speed_m2[15]), 
            .\speed_m2[16] (speed_m2[16]), .\speed_m2[17] (speed_m2[17]), 
            .\speed_m2[18] (speed_m2[18]), .\speed_m2[19] (speed_m2[19]), 
            .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(326[14:18])
    VLO i1 (.Z(GND_net));
    AVG_SPEED AVG_SPEED_M4 (.\speed_avg_m4[0] (speed_avg_m4[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m4[0] (speed_m4[0]), .\speed_avg_m4[1] (speed_avg_m4[1]), 
            .\speed_m4[1] (speed_m4[1]), .\speed_avg_m4[2] (speed_avg_m4[2]), 
            .\speed_m4[2] (speed_m4[2]), .\speed_avg_m4[3] (speed_avg_m4[3]), 
            .\speed_m4[3] (speed_m4[3]), .\speed_avg_m4[4] (speed_avg_m4[4]), 
            .\speed_m4[4] (speed_m4[4]), .\speed_avg_m4[5] (speed_avg_m4[5]), 
            .\speed_m4[5] (speed_m4[5]), .\speed_avg_m4[6] (speed_avg_m4[6]), 
            .\speed_m4[6] (speed_m4[6]), .\speed_avg_m4[7] (speed_avg_m4[7]), 
            .\speed_m4[7] (speed_m4[7]), .\speed_avg_m4[8] (speed_avg_m4[8]), 
            .\speed_m4[8] (speed_m4[8]), .\speed_avg_m4[9] (speed_avg_m4[9]), 
            .\speed_m4[9] (speed_m4[9]), .\speed_avg_m4[10] (speed_avg_m4[10]), 
            .\speed_m4[10] (speed_m4[10]), .\speed_avg_m4[11] (speed_avg_m4[11]), 
            .\speed_m4[11] (speed_m4[11]), .\speed_avg_m4[12] (speed_avg_m4[12]), 
            .\speed_m4[12] (speed_m4[12]), .\speed_avg_m4[13] (speed_avg_m4[13]), 
            .\speed_m4[13] (speed_m4[13]), .\speed_avg_m4[14] (speed_avg_m4[14]), 
            .\speed_m4[14] (speed_m4[14]), .\speed_avg_m4[15] (speed_avg_m4[15]), 
            .\speed_m4[15] (speed_m4[15]), .\speed_avg_m4[16] (speed_avg_m4[16]), 
            .\speed_m4[16] (speed_m4[16]), .\speed_avg_m4[17] (speed_avg_m4[17]), 
            .\speed_m4[17] (speed_m4[17]), .\speed_avg_m4[18] (speed_avg_m4[18]), 
            .\speed_m4[18] (speed_m4[18]), .\speed_avg_m4[19] (speed_avg_m4[19]), 
            .\speed_m4[19] (speed_m4[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(364[17:26])
    FD1P3AX start_cnt_2076__i1 (.D(n74), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i1.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i2 (.D(n73), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i2.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i3 (.D(n72), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i3.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i4 (.D(n71), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i4.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i5 (.D(n70), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i5.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i6 (.D(n69), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i6.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i7 (.D(n68), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i7.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i8 (.D(n67), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i8.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i9 (.D(n66), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i9.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i10 (.D(n65), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i10.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i11 (.D(n64), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i11.GSR = "DISABLED";
    FD1P3AX start_cnt_2076__i12 (.D(n63), .SP(clkout_c_enable_266), .CK(clkout_c), 
            .Q(start_cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i12.GSR = "DISABLED";
    FD1S3AX start_cnt_2076__i13 (.D(n10392), .CK(clkout_c), .Q(start_cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(385[18:27])
    defparam start_cnt_2076__i13.GSR = "DISABLED";
    AVG_SPEED_U9 AVG_SPEED_M3 (.\speed_avg_m3[0] (speed_avg_m3[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m3[0] (speed_m3[0]), .\speed_avg_m3[1] (speed_avg_m3[1]), 
            .\speed_m3[1] (speed_m3[1]), .\speed_avg_m3[2] (speed_avg_m3[2]), 
            .\speed_m3[2] (speed_m3[2]), .\speed_avg_m3[3] (speed_avg_m3[3]), 
            .\speed_m3[3] (speed_m3[3]), .\speed_avg_m3[4] (speed_avg_m3[4]), 
            .\speed_m3[4] (speed_m3[4]), .\speed_avg_m3[5] (speed_avg_m3[5]), 
            .\speed_m3[5] (speed_m3[5]), .\speed_avg_m3[6] (speed_avg_m3[6]), 
            .\speed_m3[6] (speed_m3[6]), .\speed_avg_m3[7] (speed_avg_m3[7]), 
            .\speed_m3[7] (speed_m3[7]), .\speed_avg_m3[8] (speed_avg_m3[8]), 
            .\speed_m3[8] (speed_m3[8]), .\speed_avg_m3[9] (speed_avg_m3[9]), 
            .\speed_m3[9] (speed_m3[9]), .\speed_avg_m3[10] (speed_avg_m3[10]), 
            .\speed_m3[10] (speed_m3[10]), .\speed_avg_m3[11] (speed_avg_m3[11]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_avg_m3[12] (speed_avg_m3[12]), 
            .\speed_m3[12] (speed_m3[12]), .\speed_avg_m3[13] (speed_avg_m3[13]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_avg_m3[14] (speed_avg_m3[14]), 
            .\speed_m3[14] (speed_m3[14]), .\speed_avg_m3[15] (speed_avg_m3[15]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_avg_m3[16] (speed_avg_m3[16]), 
            .\speed_m3[16] (speed_m3[16]), .\speed_avg_m3[17] (speed_avg_m3[17]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_avg_m3[18] (speed_avg_m3[18]), 
            .\speed_m3[18] (speed_m3[18]), .\speed_avg_m3[19] (speed_avg_m3[19]), 
            .\speed_m3[19] (speed_m3[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(361[17:26])
    AVG_SPEED_U10 AVG_SPEED_M2 (.\speed_avg_m2[0] (speed_avg_m2[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m2[0] (speed_m2[0]), .\speed_avg_m2[1] (speed_avg_m2[1]), 
            .\speed_m2[1] (speed_m2[1]), .\speed_avg_m2[2] (speed_avg_m2[2]), 
            .\speed_m2[2] (speed_m2[2]), .\speed_avg_m2[3] (speed_avg_m2[3]), 
            .\speed_m2[3] (speed_m2[3]), .\speed_avg_m2[4] (speed_avg_m2[4]), 
            .\speed_m2[4] (speed_m2[4]), .\speed_avg_m2[5] (speed_avg_m2[5]), 
            .\speed_m2[5] (speed_m2[5]), .\speed_avg_m2[6] (speed_avg_m2[6]), 
            .\speed_m2[6] (speed_m2[6]), .\speed_avg_m2[7] (speed_avg_m2[7]), 
            .\speed_m2[7] (speed_m2[7]), .\speed_avg_m2[8] (speed_avg_m2[8]), 
            .\speed_m2[8] (speed_m2[8]), .\speed_avg_m2[9] (speed_avg_m2[9]), 
            .\speed_m2[9] (speed_m2[9]), .\speed_avg_m2[10] (speed_avg_m2[10]), 
            .\speed_m2[10] (speed_m2[10]), .\speed_avg_m2[11] (speed_avg_m2[11]), 
            .\speed_m2[11] (speed_m2[11]), .\speed_avg_m2[12] (speed_avg_m2[12]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_avg_m2[13] (speed_avg_m2[13]), 
            .\speed_m2[13] (speed_m2[13]), .\speed_avg_m2[14] (speed_avg_m2[14]), 
            .\speed_m2[14] (speed_m2[14]), .\speed_avg_m2[15] (speed_avg_m2[15]), 
            .\speed_m2[15] (speed_m2[15]), .\speed_avg_m2[16] (speed_avg_m2[16]), 
            .\speed_m2[16] (speed_m2[16]), .\speed_avg_m2[17] (speed_avg_m2[17]), 
            .\speed_m2[17] (speed_m2[17]), .\speed_avg_m2[18] (speed_avg_m2[18]), 
            .\speed_m2[18] (speed_m2[18]), .\speed_avg_m2[19] (speed_avg_m2[19]), 
            .\speed_m2[19] (speed_m2[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(358[17:26])
    TSALL TSALL_INST (.TSALL(GND_net));
    AVG_SPEED_U11 AVG_SPEED_M1 (.\speed_avg_m1[0] (speed_avg_m1[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m1[0] (speed_m1[0]), .\speed_avg_m1[1] (speed_avg_m1[1]), 
            .\speed_m1[1] (speed_m1[1]), .\speed_avg_m1[2] (speed_avg_m1[2]), 
            .\speed_m1[2] (speed_m1[2]), .\speed_avg_m1[3] (speed_avg_m1[3]), 
            .\speed_m1[3] (speed_m1[3]), .\speed_avg_m1[4] (speed_avg_m1[4]), 
            .\speed_m1[4] (speed_m1[4]), .\speed_avg_m1[5] (speed_avg_m1[5]), 
            .\speed_m1[5] (speed_m1[5]), .\speed_avg_m1[6] (speed_avg_m1[6]), 
            .\speed_m1[6] (speed_m1[6]), .\speed_avg_m1[7] (speed_avg_m1[7]), 
            .\speed_m1[7] (speed_m1[7]), .\speed_avg_m1[8] (speed_avg_m1[8]), 
            .\speed_m1[8] (speed_m1[8]), .\speed_avg_m1[9] (speed_avg_m1[9]), 
            .\speed_m1[9] (speed_m1[9]), .\speed_avg_m1[10] (speed_avg_m1[10]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_avg_m1[11] (speed_avg_m1[11]), 
            .\speed_m1[11] (speed_m1[11]), .\speed_avg_m1[12] (speed_avg_m1[12]), 
            .\speed_m1[12] (speed_m1[12]), .\speed_avg_m1[13] (speed_avg_m1[13]), 
            .\speed_m1[13] (speed_m1[13]), .\speed_avg_m1[14] (speed_avg_m1[14]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_avg_m1[15] (speed_avg_m1[15]), 
            .\speed_m1[15] (speed_m1[15]), .\speed_avg_m1[16] (speed_avg_m1[16]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_avg_m1[17] (speed_avg_m1[17]), 
            .\speed_m1[17] (speed_m1[17]), .\speed_avg_m1[18] (speed_avg_m1[18]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_avg_m1[19] (speed_avg_m1[19]), 
            .\speed_m1[19] (speed_m1[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(355[17:26])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    SPI SPI_I (.GND_net(GND_net), .speed_set_m4({speed_set_m4}), .clkout_c(clkout_c), 
        .MISO_N_624(MISO_N_624), .clkout_c_enable_172(clkout_c_enable_172), 
        .enable_m1(enable_m1), .enable_m2(enable_m2), .enable_m3(enable_m3), 
        .enable_m4(enable_m4), .clkout_c_enable_173(clkout_c_enable_173), 
        .CS_c(CS_c), .SCK_c(SCK_c), .speed_set_m3({speed_set_m3}), .hallsense_m1({hallsense_m1}), 
        .dir_m1(dir_m1), .n2860(n2860), .n2896(n2896), .hallsense_m2({hallsense_m2}), 
        .dir_m2(dir_m2), .n2968(n2968), .n3004(n3004), .rst(rst), .MOSI_c(MOSI_c), 
        .hallsense_m3({hallsense_m3}), .dir_m3(dir_m3), .n3076(n3076), 
        .n3112(n3112), .n22100(n22100), .n21354(n21354), .hallsense_m4({hallsense_m4}), 
        .dir_m4(dir_m4), .n3184(n3184), .n3220(n3220), .\send_buffer[94] (send_buffer[94]), 
        .\send_buffer_95__N_346[94] (send_buffer_95__N_346[94]), .\speed_avg_m1[0] (speed_avg_m1[0]), 
        .\speed_avg_m1[8] (speed_avg_m1[8]), .\speed_avg_m1[9] (speed_avg_m1[9]), 
        .\speed_avg_m2[19] (speed_avg_m2[19]), .\speed_avg_m1[10] (speed_avg_m1[10]), 
        .\speed_avg_m1[6] (speed_avg_m1[6]), .\speed_avg_m1[7] (speed_avg_m1[7]), 
        .\speed_avg_m1[4] (speed_avg_m1[4]), .\speed_avg_m1[2] (speed_avg_m1[2]), 
        .\speed_avg_m1[1] (speed_avg_m1[1]), .\speed_avg_m1[3] (speed_avg_m1[3]), 
        .\speed_avg_m1[5] (speed_avg_m1[5]), .\speed_avg_m1[11] (speed_avg_m1[11]), 
        .\speed_avg_m1[12] (speed_avg_m1[12]), .\speed_avg_m1[13] (speed_avg_m1[13]), 
        .\speed_avg_m1[14] (speed_avg_m1[14]), .\speed_avg_m1[15] (speed_avg_m1[15]), 
        .\speed_avg_m1[16] (speed_avg_m1[16]), .\speed_avg_m1[17] (speed_avg_m1[17]), 
        .\speed_avg_m1[18] (speed_avg_m1[18]), .\speed_avg_m4[8] (speed_avg_m4[8]), 
        .\speed_avg_m4[7] (speed_avg_m4[7]), .\speed_avg_m4[10] (speed_avg_m4[10]), 
        .\speed_avg_m4[9] (speed_avg_m4[9]), .\speed_avg_m4[11] (speed_avg_m4[11]), 
        .\speed_avg_m4[12] (speed_avg_m4[12]), .\speed_avg_m4[13] (speed_avg_m4[13]), 
        .\speed_avg_m4[14] (speed_avg_m4[14]), .\speed_avg_m4[15] (speed_avg_m4[15]), 
        .\speed_avg_m4[16] (speed_avg_m4[16]), .\speed_avg_m4[17] (speed_avg_m4[17]), 
        .\speed_avg_m4[18] (speed_avg_m4[18]), .\speed_avg_m4[19] (speed_avg_m4[19]), 
        .\speed_avg_m3[0] (speed_avg_m3[0]), .\speed_avg_m3[1] (speed_avg_m3[1]), 
        .\speed_avg_m3[2] (speed_avg_m3[2]), .\speed_avg_m3[3] (speed_avg_m3[3]), 
        .\speed_avg_m3[4] (speed_avg_m3[4]), .\speed_avg_m3[5] (speed_avg_m3[5]), 
        .\speed_avg_m3[6] (speed_avg_m3[6]), .\speed_avg_m3[7] (speed_avg_m3[7]), 
        .\speed_avg_m3[8] (speed_avg_m3[8]), .\speed_avg_m3[9] (speed_avg_m3[9]), 
        .\speed_avg_m3[10] (speed_avg_m3[10]), .\speed_avg_m3[11] (speed_avg_m3[11]), 
        .speed_set_m2({speed_set_m2}), .\speed_avg_m3[12] (speed_avg_m3[12]), 
        .\speed_avg_m3[13] (speed_avg_m3[13]), .\speed_avg_m3[14] (speed_avg_m3[14]), 
        .speed_set_m1({speed_set_m1}), .\speed_avg_m3[15] (speed_avg_m3[15]), 
        .\speed_avg_m3[16] (speed_avg_m3[16]), .\speed_avg_m3[17] (speed_avg_m3[17]), 
        .\speed_avg_m3[18] (speed_avg_m3[18]), .\speed_avg_m3[19] (speed_avg_m3[19]), 
        .\speed_avg_m2[0] (speed_avg_m2[0]), .\speed_avg_m2[1] (speed_avg_m2[1]), 
        .\speed_avg_m2[2] (speed_avg_m2[2]), .\speed_avg_m2[3] (speed_avg_m2[3]), 
        .\speed_avg_m2[4] (speed_avg_m2[4]), .\speed_avg_m2[5] (speed_avg_m2[5]), 
        .\speed_avg_m2[6] (speed_avg_m2[6]), .\speed_avg_m2[7] (speed_avg_m2[7]), 
        .\speed_avg_m2[8] (speed_avg_m2[8]), .\speed_avg_m2[9] (speed_avg_m2[9]), 
        .\speed_avg_m2[10] (speed_avg_m2[10]), .\speed_avg_m2[11] (speed_avg_m2[11]), 
        .\speed_avg_m2[12] (speed_avg_m2[12]), .\speed_avg_m2[13] (speed_avg_m2[13]), 
        .\speed_avg_m2[14] (speed_avg_m2[14]), .\speed_avg_m2[15] (speed_avg_m2[15]), 
        .\speed_avg_m2[16] (speed_avg_m2[16]), .\speed_avg_m2[17] (speed_avg_m2[17]), 
        .\speed_avg_m2[18] (speed_avg_m2[18]), .\speed_avg_m4[0] (speed_avg_m4[0]), 
        .\speed_avg_m4[1] (speed_avg_m4[1]), .\speed_avg_m1[19] (speed_avg_m1[19]), 
        .\speed_avg_m4[2] (speed_avg_m4[2]), .\speed_avg_m4[3] (speed_avg_m4[3]), 
        .\speed_avg_m4[4] (speed_avg_m4[4]), .\speed_avg_m4[5] (speed_avg_m4[5]), 
        .\speed_avg_m4[6] (speed_avg_m4[6]), .n21336(n21336), .n5132(n5132), 
        .free_m4(free_m4), .n19415(n19415), .free_m3(free_m3), .n19427(n19427), 
        .free_m2(free_m2), .n19411(n19411), .free_m1(free_m1), .n19421(n19421));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(307[10:13])
    FD1S3AX rst_12_rep_409 (.D(n21309), .CK(clkout_c), .Q(n22100));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(380[3] 387[10])
    defparam rst_12_rep_409.GSR = "DISABLED";
    PWMGENERATOR_U0 PWM_I_M3 (.PWM_m3(PWM_m3), .pwm_clk(pwm_clk), .free_m3(free_m3), 
            .rst(rst), .PWMdut_m3({PWMdut_m3}), .GND_net(GND_net), .hallsense_m3({hallsense_m3}), 
            .n21363(n21363), .enable_m3(enable_m3), .n3124(n3124), .n21366(n21366), 
            .n3088(n3088));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(342[13:25])
    PWMGENERATOR_U1 PWM_I_M2 (.PWMdut_m2({PWMdut_m2}), .GND_net(GND_net), 
            .PWM_m2(PWM_m2), .pwm_clk(pwm_clk), .free_m2(free_m2), .rst(rst), 
            .hallsense_m2({hallsense_m2}), .n21369(n21369), .enable_m2(enable_m2), 
            .n3016(n3016), .n21371(n21371), .n2980(n2980));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(332[13:25])
    PWMGENERATOR_U2 PWM_I_M1 (.GND_net(GND_net), .PWM_m1(PWM_m1), .pwm_clk(pwm_clk), 
            .free_m1(free_m1), .rst(rst), .PWMdut_m1({PWMdut_m1}), .hallsense_m1({hallsense_m1}), 
            .n21373(n21373), .enable_m1(enable_m1), .n2908(n2908), .n21375(n21375), 
            .n2872(n2872));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(322[13:25])
    PWMGENERATOR PWM_I_M4 (.PWM_m4(PWM_m4), .pwm_clk(pwm_clk), .free_m4(free_m4), 
            .rst(rst), .PWMdut_m4({PWMdut_m4}), .GND_net(GND_net), .hallsense_m4({hallsense_m4}), 
            .n21358(n21358), .enable_m4(enable_m4), .n3232(n3232), .n21361(n21361), 
            .n3196(n3196));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(352[13:25])
    \PID(16000000,160000000,10000000)  PID_I (.\speed_avg_m4[5] (speed_avg_m4[5]), 
            .\speed_avg_m3[5] (speed_avg_m3[5]), .n21328(n21328), .n4322(n4322), 
            .speed_set_m2({speed_set_m2}), .speed_set_m3({speed_set_m3}), 
            .clk_N_683(clk_N_683), .n18938(n18938), .speed_set_m4({speed_set_m4}), 
            .\speed_avg_m4[18] (speed_avg_m4[18]), .\speed_avg_m3[18] (speed_avg_m3[18]), 
            .\speed_avg_m4[4] (speed_avg_m4[4]), .\speed_avg_m3[4] (speed_avg_m3[4]), 
            .\speed_avg_m3[3] (speed_avg_m3[3]), .\speed_avg_m2[3] (speed_avg_m2[3]), 
            .\speed_avg_m4[2] (speed_avg_m4[2]), .\speed_avg_m3[2] (speed_avg_m3[2]), 
            .\speed_avg_m4[1] (speed_avg_m4[1]), .\speed_avg_m3[1] (speed_avg_m3[1]), 
            .n7(n7), .GND_net(GND_net), .n4417(n4417), .n4416(n4416), 
            .\speed_avg_m4[0] (speed_avg_m4[0]), .\speed_avg_m3[0] (speed_avg_m3[0]), 
            .\speed_avg_m4[17] (speed_avg_m4[17]), .\speed_avg_m3[17] (speed_avg_m3[17]), 
            .\subOut_24__N_1177[0] (subOut_24__N_1177[0]), .speed_set_m1({speed_set_m1}), 
            .\speed_avg_m4[16] (speed_avg_m4[16]), .\speed_avg_m3[16] (speed_avg_m3[16]), 
            .\speed_avg_m4[15] (speed_avg_m4[15]), .\speed_avg_m3[15] (speed_avg_m3[15]), 
            .\speed_avg_m4[14] (speed_avg_m4[14]), .\speed_avg_m3[14] (speed_avg_m3[14]), 
            .\speed_avg_m4[13] (speed_avg_m4[13]), .\speed_avg_m3[13] (speed_avg_m3[13]), 
            .n4419(n4419), .n4418(n4418), .\speed_avg_m3[12] (speed_avg_m3[12]), 
            .\speed_avg_m2[12] (speed_avg_m2[12]), .n22100(n22100), .\speed_avg_m4[11] (speed_avg_m4[11]), 
            .\speed_avg_m3[11] (speed_avg_m3[11]), .\speed_avg_m4[10] (speed_avg_m4[10]), 
            .\speed_avg_m3[10] (speed_avg_m3[10]), .\speed_avg_m3[9] (speed_avg_m3[9]), 
            .\speed_avg_m2[9] (speed_avg_m2[9]), .n4421(n4421), .n4420(n4420), 
            .\speed_avg_m3[8] (speed_avg_m3[8]), .\speed_avg_m2[8] (speed_avg_m2[8]), 
            .n4423(n4423), .n4422(n4422), .\speed_avg_m3[7] (speed_avg_m3[7]), 
            .\speed_avg_m2[7] (speed_avg_m2[7]), .\speed_avg_m4[6] (speed_avg_m4[6]), 
            .\speed_avg_m3[6] (speed_avg_m3[6]), .n4425(n4425), .n4424(n4424), 
            .\speed_avg_m4[7] (speed_avg_m4[7]), .\speed_avg_m1[18] (speed_avg_m1[18]), 
            .\speed_avg_m2[18] (speed_avg_m2[18]), .\speed_avg_m1[17] (speed_avg_m1[17]), 
            .\speed_avg_m2[17] (speed_avg_m2[17]), .\speed_avg_m1[16] (speed_avg_m1[16]), 
            .\speed_avg_m2[16] (speed_avg_m2[16]), .\speed_avg_m1[15] (speed_avg_m1[15]), 
            .\speed_avg_m2[15] (speed_avg_m2[15]), .\speed_avg_m1[14] (speed_avg_m1[14]), 
            .\speed_avg_m2[14] (speed_avg_m2[14]), .\speed_avg_m1[13] (speed_avg_m1[13]), 
            .\speed_avg_m2[13] (speed_avg_m2[13]), .\speed_avg_m1[12] (speed_avg_m1[12]), 
            .\speed_avg_m1[11] (speed_avg_m1[11]), .\speed_avg_m2[11] (speed_avg_m2[11]), 
            .\speed_avg_m1[10] (speed_avg_m1[10]), .\speed_avg_m2[10] (speed_avg_m2[10]), 
            .\speed_avg_m1[9] (speed_avg_m1[9]), .\speed_avg_m1[8] (speed_avg_m1[8]), 
            .\speed_avg_m1[7] (speed_avg_m1[7]), .\speed_avg_m1[6] (speed_avg_m1[6]), 
            .\speed_avg_m2[6] (speed_avg_m2[6]), .\speed_avg_m1[5] (speed_avg_m1[5]), 
            .\speed_avg_m2[5] (speed_avg_m2[5]), .\speed_avg_m1[4] (speed_avg_m1[4]), 
            .\speed_avg_m2[4] (speed_avg_m2[4]), .\speed_avg_m1[3] (speed_avg_m1[3]), 
            .\speed_avg_m1[2] (speed_avg_m1[2]), .\speed_avg_m2[2] (speed_avg_m2[2]), 
            .\speed_avg_m1[1] (speed_avg_m1[1]), .\speed_avg_m2[1] (speed_avg_m2[1]), 
            .\speed_avg_m1[19] (speed_avg_m1[19]), .\speed_avg_m2[19] (speed_avg_m2[19]), 
            .n5(n5), .\speed_avg_m1[0] (speed_avg_m1[0]), .\speed_avg_m2[0] (speed_avg_m2[0]), 
            .dir_m2(dir_m2), .dir_m3(dir_m3), .dir_m1(dir_m1), .dir_m4(dir_m4), 
            .VCC_net(VCC_net), .\subOut_24__N_1177[1] (subOut_24__N_1177[1]), 
            .\subOut_24__N_1177[2] (subOut_24__N_1177[2]), .\subOut_24__N_1177[3] (subOut_24__N_1177[3]), 
            .\subOut_24__N_1177[4] (subOut_24__N_1177[4]), .\subOut_24__N_1177[5] (subOut_24__N_1177[5]), 
            .\subOut_24__N_1177[6] (subOut_24__N_1177[6]), .\subOut_24__N_1177[7] (subOut_24__N_1177[7]), 
            .\subOut_24__N_1177[8] (subOut_24__N_1177[8]), .\subOut_24__N_1177[9] (subOut_24__N_1177[9]), 
            .\subOut_24__N_1177[10] (subOut_24__N_1177[10]), .\subOut_24__N_1177[11] (subOut_24__N_1177[11]), 
            .\subOut_24__N_1177[12] (subOut_24__N_1177[12]), .\subOut_24__N_1177[13] (subOut_24__N_1177[13]), 
            .\subOut_24__N_1177[14] (subOut_24__N_1177[14]), .\subOut_24__N_1177[15] (subOut_24__N_1177[15]), 
            .\subOut_24__N_1177[16] (subOut_24__N_1177[16]), .\subOut_24__N_1177[17] (subOut_24__N_1177[17]), 
            .\subOut_24__N_1177[18] (subOut_24__N_1177[18]), .\subOut_24__N_1177[19] (subOut_24__N_1177[19]), 
            .\subOut_24__N_1177[20] (subOut_24__N_1177[20]), .\subOut_24__N_1177[21] (subOut_24__N_1177[21]), 
            .\subOut_24__N_1177[24] (subOut_24__N_1177[24]), .n4427(n4427), 
            .n4426(n4426), .n4429(n4429), .n4428(n4428), .n4431(n4431), 
            .n4430(n4430), .n4433(n4433), .n4432(n4432), .n20284(n20284), 
            .n4435(n4435), .n4434(n4434), .n4436(n4436), .n4440(n4440), 
            .n4442(n4442), .n4441(n4441), .n4444(n4444), .n4443(n4443), 
            .n4446(n4446), .n4445(n4445), .PWMdut_m4({PWMdut_m4}), .PWMdut_m3({PWMdut_m3}), 
            .PWMdut_m2({PWMdut_m2}), .n4448(n4448), .n4447(n4447), .n4450(n4450), 
            .n4449(n4449), .PWMdut_m1({PWMdut_m1}), .n4452(n4452), .n4451(n4451), 
            .n4454(n4454), .n4453(n4453), .n4456(n4456), .n4455(n4455), 
            .\speed_avg_m4[3] (speed_avg_m4[3]), .n4458(n4458), .n4457(n4457), 
            .n4460(n4460), .n4459(n4459), .n4461(n4461), .\speed_avg_m4[12] (speed_avg_m4[12]), 
            .\speed_avg_m4[9] (speed_avg_m4[9]), .\speed_avg_m4[8] (speed_avg_m4[8]), 
            .n4415(n4415), .n4414(n4414));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(311[10:13])
    HALL_U5 HALL_I_M1 (.clk_1mhz(clk_1mhz), .n22097(n22097), .\speed_m1[0] (speed_m1[0]), 
            .hallsense_m1({hallsense_m1}), .rst(rst), .clkout_c_enable_173(clkout_c_enable_173), 
            .H_A_m1_c(H_A_m1_c), .H_B_m1_c(H_B_m1_c), .H_C_m1_c(H_C_m1_c), 
            .\speed_m1[1] (speed_m1[1]), .\speed_m1[2] (speed_m1[2]), .\speed_m1[3] (speed_m1[3]), 
            .\speed_m1[4] (speed_m1[4]), .\speed_m1[5] (speed_m1[5]), .\speed_m1[6] (speed_m1[6]), 
            .\speed_m1[7] (speed_m1[7]), .\speed_m1[8] (speed_m1[8]), .\speed_m1[9] (speed_m1[9]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_m1[11] (speed_m1[11]), 
            .\speed_m1[12] (speed_m1[12]), .\speed_m1[13] (speed_m1[13]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_m1[15] (speed_m1[15]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_m1[17] (speed_m1[17]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_m1[19] (speed_m1[19]), 
            .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(316[14:18])
    HALL_U3 HALL_I_M3 (.\speed_m3[0] (speed_m3[0]), .clk_1mhz(clk_1mhz), 
            .hallsense_m3({hallsense_m3}), .clkout_c_enable_173(clkout_c_enable_173), 
            .H_A_m3_c(H_A_m3_c), .H_B_m3_c(H_B_m3_c), .H_C_m3_c(H_C_m3_c), 
            .rst(rst), .\speed_m3[1] (speed_m3[1]), .\speed_m3[2] (speed_m3[2]), 
            .\speed_m3[3] (speed_m3[3]), .\speed_m3[4] (speed_m3[4]), .\speed_m3[5] (speed_m3[5]), 
            .\speed_m3[6] (speed_m3[6]), .\speed_m3[7] (speed_m3[7]), .\speed_m3[8] (speed_m3[8]), 
            .\speed_m3[9] (speed_m3[9]), .\speed_m3[10] (speed_m3[10]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_m3[12] (speed_m3[12]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_m3[14] (speed_m3[14]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_m3[16] (speed_m3[16]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_m3[18] (speed_m3[18]), 
            .\speed_m3[19] (speed_m3[19]), .GND_net(GND_net), .n22097(n22097));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(336[14:18])
    HALL HALL_I_M4 (.clk_1mhz(clk_1mhz), .\speed_m4[0] (speed_m4[0]), .hallsense_m4({hallsense_m4}), 
         .clkout_c_enable_172(clkout_c_enable_172), .clkout_c_enable_173(clkout_c_enable_173), 
         .HALL_A_OUT_c_c(HALL_A_OUT_c_c), .HALL_B_OUT_c_c(HALL_B_OUT_c_c), 
         .rst(rst), .HALL_C_OUT_c_c(HALL_C_OUT_c_c), .\speed_m4[1] (speed_m4[1]), 
         .\speed_m4[2] (speed_m4[2]), .\speed_m4[3] (speed_m4[3]), .\speed_m4[4] (speed_m4[4]), 
         .\speed_m4[5] (speed_m4[5]), .\speed_m4[6] (speed_m4[6]), .\speed_m4[7] (speed_m4[7]), 
         .\speed_m4[8] (speed_m4[8]), .\speed_m4[9] (speed_m4[9]), .\speed_m4[10] (speed_m4[10]), 
         .\speed_m4[11] (speed_m4[11]), .\speed_m4[12] (speed_m4[12]), .\speed_m4[13] (speed_m4[13]), 
         .\speed_m4[14] (speed_m4[14]), .\speed_m4[15] (speed_m4[15]), .\speed_m4[16] (speed_m4[16]), 
         .\speed_m4[17] (speed_m4[17]), .\speed_m4[18] (speed_m4[18]), .\speed_m4[19] (speed_m4[19]), 
         .GND_net(GND_net), .n22097(n22097));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(346[14:18])
    
endmodule
//
// Verilog Description of module COMMUTATION_U6
//

module COMMUTATION_U6 (MB_m3_c_0, clkout_c, MC_m3_c_0, MA_m3_c_0, LED3_c, 
            enable_m3, n3076, n21366, PWM_m3, n3112, n21363, n19427, 
            n21362, free_m3, MA_m3_c_1, n3170, MC_m3_c_1, n3124, 
            MB_m3_c_1, n3088);
    output MB_m3_c_0;
    input clkout_c;
    output MC_m3_c_0;
    output MA_m3_c_0;
    output LED3_c;
    input enable_m3;
    input n3076;
    input n21366;
    input PWM_m3;
    input n3112;
    input n21363;
    input n19427;
    input n21362;
    input free_m3;
    output MA_m3_c_1;
    input n3170;
    output MC_m3_c_1;
    input n3124;
    output MB_m3_c_1;
    input n3088;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1957, n18518, n18517, n19428, n14093;
    
    FD1S3IX MospairB_i1 (.D(n18518), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MB_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18517), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MC_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19428), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MA_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14093), .CK(clkout_c), .PD(led1_N_1957), .Q(LED3_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10618_1_lut (.A(enable_m3), .Z(led1_N_1957)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10618_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3076), .B(n21366), .C(PWM_m3), .Z(n18518)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_176 (.A(n3112), .B(n21363), .C(PWM_m3), .Z(n18517)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_176.init = 16'hbfbf;
    LUT4 i17130_3_lut (.A(n19427), .B(PWM_m3), .C(n21362), .Z(n19428)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17130_3_lut.init = 16'hbfbf;
    LUT4 i11521_2_lut (.A(free_m3), .B(LED3_c), .Z(n14093)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11521_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n3170), .CK(clkout_c), .CD(n19427), .Q(MA_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3112), .CK(clkout_c), .CD(n3124), .Q(MC_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3076), .CK(clkout_c), .CD(n3088), .Q(MB_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION_U7
//

module COMMUTATION_U7 (MB_m2_c_0, clkout_c, MC_m2_c_0, MA_m2_c_0, LED2_c, 
            enable_m2, n2968, n21371, PWM_m2, n3004, n21369, n19411, 
            n21368, free_m2, MA_m2_c_1, n3062, MC_m2_c_1, n3016, 
            MB_m2_c_1, n2980);
    output MB_m2_c_0;
    input clkout_c;
    output MC_m2_c_0;
    output MA_m2_c_0;
    output LED2_c;
    input enable_m2;
    input n2968;
    input n21371;
    input PWM_m2;
    input n3004;
    input n21369;
    input n19411;
    input n21368;
    input free_m2;
    output MA_m2_c_1;
    input n3062;
    output MC_m2_c_1;
    input n3016;
    output MB_m2_c_1;
    input n2980;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1957, n18520, n18519, n19412, n14095;
    
    FD1S3IX MospairB_i1 (.D(n18520), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MB_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18519), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MC_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19412), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MA_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14095), .CK(clkout_c), .PD(led1_N_1957), .Q(LED2_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10617_1_lut (.A(enable_m2), .Z(led1_N_1957)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10617_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2968), .B(n21371), .C(PWM_m2), .Z(n18520)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_175 (.A(n3004), .B(n21369), .C(PWM_m2), .Z(n18519)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_175.init = 16'hbfbf;
    LUT4 i17133_3_lut (.A(n19411), .B(PWM_m2), .C(n21368), .Z(n19412)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17133_3_lut.init = 16'hbfbf;
    LUT4 i11523_2_lut (.A(free_m2), .B(LED2_c), .Z(n14095)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11523_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n3062), .CK(clkout_c), .CD(n19411), .Q(MA_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3004), .CK(clkout_c), .CD(n3016), .Q(MC_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2968), .CK(clkout_c), .CD(n2980), .Q(MB_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=329, LSE_RLINE=329 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION_U8
//

module COMMUTATION_U8 (MB_m1_c_0, clkout_c, MC_m1_c_0, MA_m1_c_0, LED1_c, 
            enable_m1, n2860, n21375, PWM_m1, n2896, n21373, n19421, 
            n21372, free_m1, MA_m1_c_1, n2954, MC_m1_c_1, n2908, 
            MB_m1_c_1, n2872);
    output MB_m1_c_0;
    input clkout_c;
    output MC_m1_c_0;
    output MA_m1_c_0;
    output LED1_c;
    input enable_m1;
    input n2860;
    input n21375;
    input PWM_m1;
    input n2896;
    input n21373;
    input n19421;
    input n21372;
    input free_m1;
    output MA_m1_c_1;
    input n2954;
    output MC_m1_c_1;
    input n2908;
    output MB_m1_c_1;
    input n2872;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1957, n18522, n18521, n19422, n14097;
    
    FD1S3IX MospairB_i1 (.D(n18522), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MB_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18521), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MC_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19422), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MA_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14097), .CK(clkout_c), .PD(led1_N_1957), .Q(LED1_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10616_1_lut (.A(enable_m1), .Z(led1_N_1957)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10616_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n2860), .B(n21375), .C(PWM_m1), .Z(n18522)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_174 (.A(n2896), .B(n21373), .C(PWM_m1), .Z(n18521)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_174.init = 16'hbfbf;
    LUT4 i17136_3_lut (.A(n19421), .B(PWM_m1), .C(n21372), .Z(n19422)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17136_3_lut.init = 16'hbfbf;
    LUT4 i11525_2_lut (.A(free_m1), .B(LED1_c), .Z(n14097)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11525_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n2954), .CK(clkout_c), .CD(n19421), .Q(MA_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n2896), .CK(clkout_c), .CD(n2908), .Q(MC_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n2860), .CK(clkout_c), .CD(n2872), .Q(MB_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=319, LSE_RLINE=319 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module CLKDIV
//

module CLKDIV (clkout_c, clk_1mhz, pwm_clk, GND_net, clk_N_683);
    input clkout_c;
    output clk_1mhz;
    output pwm_clk;
    input GND_net;
    output clk_N_683;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    wire pi_clk /* synthesis is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(89[9:15])
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    wire [4:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(41[8:13])
    
    wire n19716, n14136, pi_buf, n14135, pi_buf_N_69, mhz_buf, mhz_buf_N_68, 
        n19710;
    wire [11:0]cntpi;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(42[8:13])
    
    wire n19780, pwm_buf, pwm_buf_N_67, n21348;
    wire [4:0]n25;
    wire [8:0]n41;
    
    wire n18173, n18172, n18171, n18170;
    
    LUT4 i17108_4_lut (.A(count[2]), .B(count[0]), .C(count[3]), .D(n19716), 
         .Z(n14136)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(61[5:15])
    defparam i17108_4_lut.init = 16'h0400;
    LUT4 i16328_2_lut (.A(count[4]), .B(count[1]), .Z(n19716)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16328_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(pi_buf), .B(n14135), .Z(pi_buf_N_69)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    FD1S3AX mhz_buf_29 (.D(mhz_buf_N_68), .CK(clkout_c), .Q(mhz_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam mhz_buf_29.GSR = "DISABLED";
    LUT4 i17105_4_lut (.A(n19710), .B(cntpi[2]), .C(n19780), .D(cntpi[7]), 
         .Z(n14135)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(66[5:16])
    defparam i17105_4_lut.init = 16'h0020;
    FD1S3AX pi_buf_30 (.D(pi_buf_N_69), .CK(clkout_c), .Q(pi_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pi_buf_30.GSR = "DISABLED";
    FD1S3AX pwm_buf_32 (.D(pwm_buf_N_67), .CK(clkout_c), .Q(pwm_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pwm_buf_32.GSR = "DISABLED";
    FD1S3AX clk_1mhz_33 (.D(mhz_buf), .CK(clkout_c), .Q(clk_1mhz)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam clk_1mhz_33.GSR = "DISABLED";
    FD1S3AX pwm_clk_34 (.D(pwm_buf), .CK(clkout_c), .Q(pwm_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pwm_clk_34.GSR = "DISABLED";
    FD1S3AX pi_clk_35 (.D(pi_buf), .CK(clkout_c), .Q(pi_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=302, LSE_RLINE=302 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pi_clk_35.GSR = "DISABLED";
    LUT4 i16322_3_lut (.A(cntpi[5]), .B(cntpi[3]), .C(cntpi[6]), .Z(n19710)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16322_3_lut.init = 16'h8080;
    LUT4 i16391_4_lut (.A(cntpi[1]), .B(cntpi[0]), .C(cntpi[8]), .D(cntpi[4]), 
         .Z(n19780)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16391_4_lut.init = 16'h8000;
    LUT4 pwm_buf_I_0_1_lut (.A(pwm_buf), .Z(pwm_buf_N_67)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(73[14:25])
    defparam pwm_buf_I_0_1_lut.init = 16'h5555;
    LUT4 i15045_3_lut_4_lut (.A(count[2]), .B(n21348), .C(count[3]), .D(count[4]), 
         .Z(n25[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15045_3_lut_4_lut.init = 16'h7f80;
    FD1S3IX cntpi_2078_2079__i2 (.D(n41[1]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i2.GSR = "DISABLED";
    LUT4 i15027_2_lut_rep_367 (.A(count[1]), .B(count[0]), .Z(n21348)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15027_2_lut_rep_367.init = 16'h8888;
    LUT4 i15031_2_lut_3_lut (.A(count[1]), .B(count[0]), .C(count[2]), 
         .Z(n25[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15031_2_lut_3_lut.init = 16'h7878;
    LUT4 i15038_2_lut_3_lut_4_lut (.A(count[1]), .B(count[0]), .C(count[3]), 
         .D(count[2]), .Z(n25[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15038_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D cntpi_2078_2079_add_4_9 (.A0(cntpi[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18173), .S0(n41[7]), .S1(n41[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079_add_4_9.INIT0 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_9.INIT1 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_9.INJECT1_0 = "NO";
    defparam cntpi_2078_2079_add_4_9.INJECT1_1 = "NO";
    CCU2D cntpi_2078_2079_add_4_7 (.A0(cntpi[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18172), .COUT(n18173), .S0(n41[5]), .S1(n41[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079_add_4_7.INIT0 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_7.INIT1 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_7.INJECT1_0 = "NO";
    defparam cntpi_2078_2079_add_4_7.INJECT1_1 = "NO";
    CCU2D cntpi_2078_2079_add_4_5 (.A0(cntpi[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18171), .COUT(n18172), .S0(n41[3]), .S1(n41[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079_add_4_5.INIT0 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_5.INIT1 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_5.INJECT1_0 = "NO";
    defparam cntpi_2078_2079_add_4_5.INJECT1_1 = "NO";
    CCU2D cntpi_2078_2079_add_4_3 (.A0(cntpi[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18170), .COUT(n18171), .S0(n41[1]), .S1(n41[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079_add_4_3.INIT0 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_3.INIT1 = 16'hfaaa;
    defparam cntpi_2078_2079_add_4_3.INJECT1_0 = "NO";
    defparam cntpi_2078_2079_add_4_3.INJECT1_1 = "NO";
    CCU2D cntpi_2078_2079_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18170), .S1(n41[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079_add_4_1.INIT0 = 16'hF000;
    defparam cntpi_2078_2079_add_4_1.INIT1 = 16'h0555;
    defparam cntpi_2078_2079_add_4_1.INJECT1_0 = "NO";
    defparam cntpi_2078_2079_add_4_1.INJECT1_1 = "NO";
    FD1S3IX count_2077__i0 (.D(n25[0]), .CK(clkout_c), .CD(n14136), .Q(count[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2077__i0.GSR = "DISABLED";
    FD1S3IX cntpi_2078_2079__i1 (.D(n41[0]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i1.GSR = "DISABLED";
    LUT4 i15022_1_lut (.A(count[0]), .Z(n25[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15022_1_lut.init = 16'h5555;
    LUT4 i15024_2_lut (.A(count[1]), .B(count[0]), .Z(n25[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15024_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_173 (.A(mhz_buf), .B(n14136), .Z(mhz_buf_N_68)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_173.init = 16'h6666;
    INV i17492 (.A(pi_clk), .Z(clk_N_683));
    FD1S3IX cntpi_2078_2079__i3 (.D(n41[2]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i3.GSR = "DISABLED";
    FD1S3IX cntpi_2078_2079__i4 (.D(n41[3]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i4.GSR = "DISABLED";
    FD1S3IX cntpi_2078_2079__i5 (.D(n41[4]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i5.GSR = "DISABLED";
    FD1S3IX cntpi_2078_2079__i6 (.D(n41[5]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i6.GSR = "DISABLED";
    FD1S3IX cntpi_2078_2079__i7 (.D(n41[6]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i7.GSR = "DISABLED";
    FD1S3IX cntpi_2078_2079__i8 (.D(n41[7]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i8.GSR = "DISABLED";
    FD1S3IX cntpi_2078_2079__i9 (.D(n41[8]), .CK(clkout_c), .CD(n14135), 
            .Q(cntpi[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2078_2079__i9.GSR = "DISABLED";
    FD1S3IX count_2077__i1 (.D(n25[1]), .CK(clkout_c), .CD(n14136), .Q(count[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2077__i1.GSR = "DISABLED";
    FD1S3IX count_2077__i2 (.D(n25[2]), .CK(clkout_c), .CD(n14136), .Q(count[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2077__i2.GSR = "DISABLED";
    FD1S3IX count_2077__i3 (.D(n25[3]), .CK(clkout_c), .CD(n14136), .Q(count[3]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2077__i3.GSR = "DISABLED";
    FD1S3IX count_2077__i4 (.D(n25[4]), .CK(clkout_c), .CD(n14136), .Q(count[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2077__i4.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION
//

module COMMUTATION (MB_m4_c_0, clkout_c, MC_m4_c_0, MA_m4_c_0, LED4_c, 
            enable_m4, n3184, n21361, PWM_m4, n3220, n21358, n19415, 
            n21357, free_m4, MA_m4_c_1, n3278, MC_m4_c_1, n3232, 
            MB_m4_c_1, n3196);
    output MB_m4_c_0;
    input clkout_c;
    output MC_m4_c_0;
    output MA_m4_c_0;
    output LED4_c;
    input enable_m4;
    input n3184;
    input n21361;
    input PWM_m4;
    input n3220;
    input n21358;
    input n19415;
    input n21357;
    input free_m4;
    output MA_m4_c_1;
    input n3278;
    output MC_m4_c_1;
    input n3232;
    output MB_m4_c_1;
    input n3196;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire led1_N_1957, n18516, n18515, n19416, n14091;
    
    FD1S3IX MospairB_i1 (.D(n18516), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MB_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i1 (.D(n18515), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MC_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i1.GSR = "DISABLED";
    FD1S3IX MospairA_i1 (.D(n19416), .CK(clkout_c), .CD(led1_N_1957), 
            .Q(MA_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3JX led1_46 (.D(n14091), .CK(clkout_c), .PD(led1_N_1957), .Q(LED4_c)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam led1_46.GSR = "DISABLED";
    LUT4 i10621_1_lut (.A(enable_m4), .Z(led1_N_1957)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i10621_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n3184), .B(n21361), .C(PWM_m4), .Z(n18516)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_adj_172 (.A(n3220), .B(n21358), .C(PWM_m4), .Z(n18515)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(71[3] 192[10])
    defparam i2_3_lut_adj_172.init = 16'hbfbf;
    LUT4 i17127_3_lut (.A(n19415), .B(PWM_m4), .C(n21357), .Z(n19416)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i17127_3_lut.init = 16'hbfbf;
    LUT4 i11519_2_lut (.A(free_m4), .B(LED4_c), .Z(n14091)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam i11519_2_lut.init = 16'h8888;
    FD1S3IX MospairA_i2 (.D(n3278), .CK(clkout_c), .CD(n19415), .Q(MA_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairA_i2.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n3220), .CK(clkout_c), .CD(n3232), .Q(MC_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n3184), .CK(clkout_c), .CD(n3196), .Q(MB_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=349, LSE_RLINE=349 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[2] 193[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module HALL_U4
//

module HALL_U4 (clk_1mhz, n22097, \speed_m2[0] , hallsense_m2, clkout_c_enable_173, 
            H_C_m2_c, rst, H_A_m2_c, H_B_m2_c, \speed_m2[1] , \speed_m2[2] , 
            \speed_m2[3] , \speed_m2[4] , \speed_m2[5] , \speed_m2[6] , 
            \speed_m2[7] , \speed_m2[8] , \speed_m2[9] , \speed_m2[10] , 
            \speed_m2[11] , \speed_m2[12] , \speed_m2[13] , \speed_m2[14] , 
            \speed_m2[15] , \speed_m2[16] , \speed_m2[17] , \speed_m2[18] , 
            \speed_m2[19] , GND_net);
    input clk_1mhz;
    input n22097;
    output \speed_m2[0] ;
    output [2:0]hallsense_m2;
    input clkout_c_enable_173;
    input H_C_m2_c;
    input rst;
    input H_A_m2_c;
    input H_B_m2_c;
    output \speed_m2[1] ;
    output \speed_m2[2] ;
    output \speed_m2[3] ;
    output \speed_m2[4] ;
    output \speed_m2[5] ;
    output \speed_m2[6] ;
    output \speed_m2[7] ;
    output \speed_m2[8] ;
    output \speed_m2[9] ;
    output \speed_m2[10] ;
    output \speed_m2[11] ;
    output \speed_m2[12] ;
    output \speed_m2[13] ;
    output \speed_m2[14] ;
    output \speed_m2[15] ;
    output \speed_m2[16] ;
    output \speed_m2[17] ;
    output \speed_m2[18] ;
    output \speed_m2[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire stable_counting, clk_1mhz_enable_4, n14371;
    wire [19:0]speedt_19__N_1853;
    
    wire hall3_lat;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4551;
    wire [19:0]count_19__N_1873;
    
    wire hall3_old;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_177;
    wire [6:0]n63;
    
    wire n19505, n4, stable_counting_N_1935;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n15733, n21345, n21305, n4_adj_2234, n21329, n13, n19812, 
        n11431, n19784, n19730, n19726, n19572, n19394, n11429, 
        hall1_old, hall1_lat, hall2_old, hall2_lat, n21384, n18092, 
        n18091, n18090, n18089, n18088, n18087, n18086, n18085, 
        n18084, n18083, n21327, n18693, n19632, n21, n26, n22, 
        n19746, n24, n18;
    
    FD1P3IX stable_counting_62 (.D(n22097), .SP(clk_1mhz_enable_4), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1853[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_19__N_1873[0]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX speedt_i0_i0 (.D(count_19__N_1873[0]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n63[2]), .B(n19505), .C(n63[4]), .D(n4), .Z(stable_counting_N_1935)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut.init = 16'h0004;
    LUT4 i2410_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2410_2_lut.init = 16'h6666;
    LUT4 i13183_2_lut (.A(count[0]), .B(count[10]), .Z(n15733)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13183_2_lut.init = 16'h8888;
    FD1P3AX hall3_lat_59 (.D(H_C_m2_c), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    LUT4 i2438_2_lut_rep_324_3_lut_4_lut (.A(stable_count[3]), .B(n21345), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21305)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2438_2_lut_rep_324_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2_3_lut_rep_348 (.A(hall3_old), .B(n4_adj_2234), .C(hall3_lat), 
         .Z(n21329)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_348.init = 16'hdede;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4_adj_2234), .C(hall3_lat), 
         .D(n63[1]), .Z(n19505)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 i7_4_lut (.A(n13), .B(n15733), .C(count[2]), .D(n19812), .Z(n11431)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i7_4_lut.init = 16'h0080;
    LUT4 i5_4_lut (.A(count[9]), .B(count[3]), .C(count[8]), .D(count[13]), 
         .Z(n13)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i16420_4_lut (.A(count[18]), .B(n19784), .C(n19730), .D(count[1]), 
         .Z(n19812)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16420_4_lut.init = 16'hfffe;
    LUT4 i16394_4_lut (.A(count[17]), .B(n19726), .C(n19572), .D(count[12]), 
         .Z(n19784)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16394_4_lut.init = 16'hfffe;
    LUT4 i16342_3_lut (.A(count[15]), .B(count[5]), .C(count[16]), .Z(n19730)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16342_3_lut.init = 16'hfefe;
    LUT4 i16338_4_lut (.A(count[11]), .B(count[7]), .C(count[4]), .D(count[6]), 
         .Z(n19726)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16338_4_lut.init = 16'hfffe;
    LUT4 i16188_2_lut (.A(count[19]), .B(count[14]), .Z(n19572)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16188_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(n63[4]), .B(stable_count[0]), .C(n19394), .D(n19505), 
         .Z(n11429)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(rst), .CK(clk_1mhz), .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(rst), .CK(clk_1mhz), .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m2_c), .SP(rst), .CK(clk_1mhz), .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m2_c), .SP(rst), .CK(clk_1mhz), .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    LUT4 i2242_2_lut (.A(stable_counting), .B(stable_counting_N_1935), .Z(n4551)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2242_2_lut.init = 16'h8888;
    FD1P3AX speed__i2 (.D(speedt_19__N_1853[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1853[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1853[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1853[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1853[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1853[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1853[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1853[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1853[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1853[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1853[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1853[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1853[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1853[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1853[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1853[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1853[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1853[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1853[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(count_19__N_1873[1]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_1873[2]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_1873[3]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_1873[4]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_1873[5]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_1873[6]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_1873[7]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_1873[8]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_1873[9]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_1873[10]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_1873[11]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_1873[12]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_1873[13]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_1873[14]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_1873[15]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_1873[16]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_1873[17]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_1873[18]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_1873[19]), .CK(clk_1mhz), .CD(n4551), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_1873[1]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_1873[2]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_1873[3]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_1873[4]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_1873[5]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_1873[6]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_1873[7]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_1873[8]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_1873[9]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_1873[10]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_1873[11]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_1873[12]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_1873[13]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_1873[14]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_1873[15]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_1873[16]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_1873[17]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_1873[18]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_1873[19]), .SP(clk_1mhz_enable_177), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    LUT4 i2431_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21384), .C(stable_count[4]), 
         .D(stable_count[3]), .Z(n63[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2431_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i11518_4_lut (.A(n11431), .B(n11429), .C(stable_counting), .D(stable_counting_N_1935), 
         .Z(clk_1mhz_enable_177)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11518_4_lut.init = 16'hcaea;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[0]), 
         .D(speedt[0]), .Z(speedt_19__N_1853[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[1]), 
         .D(speedt[1]), .Z(speedt_19__N_1853[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[2]), 
         .D(speedt[2]), .Z(speedt_19__N_1853[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[3]), 
         .D(speedt[3]), .Z(speedt_19__N_1853[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[4]), 
         .D(speedt[4]), .Z(speedt_19__N_1853[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[5]), 
         .D(speedt[5]), .Z(speedt_19__N_1853[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[6]), 
         .D(speedt[6]), .Z(speedt_19__N_1853[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[7]), 
         .D(speedt[7]), .Z(speedt_19__N_1853[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[8]), 
         .D(speedt[8]), .Z(speedt_19__N_1853[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[9]), 
         .D(speedt[9]), .Z(speedt_19__N_1853[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2412_2_lut_rep_403 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21384)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2412_2_lut_rep_403.init = 16'h8888;
    LUT4 i2417_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2417_2_lut_3_lut.init = 16'h7878;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18092), 
          .S0(count_19__N_1873[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18091), .COUT(n18092), .S0(count_19__N_1873[17]), .S1(count_19__N_1873[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18090), .COUT(n18091), .S0(count_19__N_1873[15]), .S1(count_19__N_1873[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[10]), 
         .D(speedt[10]), .Z(speedt_19__N_1853[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[11]), 
         .D(speedt[11]), .Z(speedt_19__N_1853[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18089), .COUT(n18090), .S0(count_19__N_1873[13]), .S1(count_19__N_1873[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[12]), 
         .D(speedt[12]), .Z(speedt_19__N_1853[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[13]), 
         .D(speedt[13]), .Z(speedt_19__N_1853[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[14]), 
         .D(speedt[14]), .Z(speedt_19__N_1853[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[15]), 
         .D(speedt[15]), .Z(speedt_19__N_1853[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18088), .COUT(n18089), .S0(count_19__N_1873[11]), .S1(count_19__N_1873[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[16]), 
         .D(speedt[16]), .Z(speedt_19__N_1853[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[17]), 
         .D(speedt[17]), .Z(speedt_19__N_1853[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[18]), 
         .D(speedt[18]), .Z(speedt_19__N_1853[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11431), .B(n11429), .C(count_19__N_1873[19]), 
         .D(speedt[19]), .Z(speedt_19__N_1853[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18087), .COUT(n18088), .S0(count_19__N_1873[9]), .S1(count_19__N_1873[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18086), 
          .COUT(n18087), .S0(count_19__N_1873[7]), .S1(count_19__N_1873[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18085), 
          .COUT(n18086), .S0(count_19__N_1873[5]), .S1(count_19__N_1873[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18084), 
          .COUT(n18085), .S0(count_19__N_1873[3]), .S1(count_19__N_1873[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18083), 
          .COUT(n18084), .S0(count_19__N_1873[1]), .S1(count_19__N_1873[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18083), 
          .S1(count_19__N_1873[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21305), .SP(stable_counting), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n63[4]), .SP(stable_counting), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_167 (.A(n63[6]), .B(n63[3]), .C(n21305), .D(stable_count[0]), 
         .Z(n4)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_167.init = 16'hfeff;
    LUT4 i1_2_lut_4_lut_adj_168 (.A(n63[6]), .B(n63[3]), .C(n21305), .D(n63[2]), 
         .Z(n19394)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_168.init = 16'hfffe;
    LUT4 i2419_2_lut_rep_364_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21345)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2419_2_lut_rep_364_3_lut.init = 16'h8080;
    LUT4 i2426_2_lut_rep_346_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21327)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2426_2_lut_rep_346_3_lut_4_lut.init = 16'h8000;
    LUT4 i2424_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2424_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14371), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=326, LSE_RLINE=326 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    LUT4 i2408_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2408_1_lut.init = 16'h5555;
    LUT4 i17084_4_lut (.A(n18693), .B(n19632), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_4)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17084_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_169 (.A(n21), .B(n15733), .C(n26), .D(n22), .Z(n18693)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i1_4_lut_adj_169.init = 16'hfffb;
    LUT4 i16247_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19632)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16247_4_lut.init = 16'h7bde;
    LUT4 i7_4_lut_adj_170 (.A(count[11]), .B(count[8]), .C(n19746), .D(count[13]), 
         .Z(n21)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i7_4_lut_adj_170.init = 16'hbfff;
    LUT4 i12_4_lut (.A(count[14]), .B(n24), .C(n18), .D(count[17]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[7]), .B(count[16]), .C(count[18]), .D(count[6]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i16357_3_lut (.A(count[2]), .B(count[3]), .C(count[9]), .Z(n19746)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16357_3_lut.init = 16'h8080;
    LUT4 i10_4_lut (.A(count[19]), .B(count[12]), .C(count[4]), .D(count[15]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[1]), .B(count[5]), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i16369_3_lut (.A(n21329), .B(stable_counting), .C(stable_counting_N_1935), 
         .Z(n14371)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16369_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_171 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4_adj_2234)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_171.init = 16'h7bde;
    LUT4 i2445_3_lut_4_lut (.A(stable_count[4]), .B(n21327), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2445_3_lut_4_lut.init = 16'h7f80;
    
endmodule
//
// Verilog Description of module AVG_SPEED
//

module AVG_SPEED (\speed_avg_m4[0] , clk_1mhz, \speed_m4[0] , \speed_avg_m4[1] , 
            \speed_m4[1] , \speed_avg_m4[2] , \speed_m4[2] , \speed_avg_m4[3] , 
            \speed_m4[3] , \speed_avg_m4[4] , \speed_m4[4] , \speed_avg_m4[5] , 
            \speed_m4[5] , \speed_avg_m4[6] , \speed_m4[6] , \speed_avg_m4[7] , 
            \speed_m4[7] , \speed_avg_m4[8] , \speed_m4[8] , \speed_avg_m4[9] , 
            \speed_m4[9] , \speed_avg_m4[10] , \speed_m4[10] , \speed_avg_m4[11] , 
            \speed_m4[11] , \speed_avg_m4[12] , \speed_m4[12] , \speed_avg_m4[13] , 
            \speed_m4[13] , \speed_avg_m4[14] , \speed_m4[14] , \speed_avg_m4[15] , 
            \speed_m4[15] , \speed_avg_m4[16] , \speed_m4[16] , \speed_avg_m4[17] , 
            \speed_m4[17] , \speed_avg_m4[18] , \speed_m4[18] , \speed_avg_m4[19] , 
            \speed_m4[19] , GND_net);
    output \speed_avg_m4[0] ;
    input clk_1mhz;
    input \speed_m4[0] ;
    output \speed_avg_m4[1] ;
    input \speed_m4[1] ;
    output \speed_avg_m4[2] ;
    input \speed_m4[2] ;
    output \speed_avg_m4[3] ;
    input \speed_m4[3] ;
    output \speed_avg_m4[4] ;
    input \speed_m4[4] ;
    output \speed_avg_m4[5] ;
    input \speed_m4[5] ;
    output \speed_avg_m4[6] ;
    input \speed_m4[6] ;
    output \speed_avg_m4[7] ;
    input \speed_m4[7] ;
    output \speed_avg_m4[8] ;
    input \speed_m4[8] ;
    output \speed_avg_m4[9] ;
    input \speed_m4[9] ;
    output \speed_avg_m4[10] ;
    input \speed_m4[10] ;
    output \speed_avg_m4[11] ;
    input \speed_m4[11] ;
    output \speed_avg_m4[12] ;
    input \speed_m4[12] ;
    output \speed_avg_m4[13] ;
    input \speed_m4[13] ;
    output \speed_avg_m4[14] ;
    input \speed_m4[14] ;
    output \speed_avg_m4[15] ;
    input \speed_m4[15] ;
    output \speed_avg_m4[16] ;
    input \speed_m4[16] ;
    output \speed_avg_m4[17] ;
    input \speed_m4[17] ;
    output \speed_avg_m4[18] ;
    input \speed_m4[18] ;
    output \speed_avg_m4[19] ;
    input \speed_m4[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_139;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n19742, n6, n18184, n18183, n18182;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m4[0] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2093__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_139), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093__i0.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m4[1] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m4[2] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m4[3] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m4[4] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m4[5] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m4[6] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m4[7] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m4[8] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m4[9] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m4[10] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m4[11] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m4[12] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m4[13] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m4[14] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m4[15] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m4[16] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m4[17] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m4[18] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m4[19] ), .SP(clk_1mhz_enable_139), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    LUT4 i17184_4_lut (.A(clk_cnt[0]), .B(n19742), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_139)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17184_4_lut.init = 16'h0004;
    LUT4 i16353_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n19742)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16353_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    CCU2D clk_cnt_2093_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18184), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2093_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2093_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2093_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2093_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18183), .COUT(n18184), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2093_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2093_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2093_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2093_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18182), .COUT(n18183), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2093_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2093_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2093_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2093_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18182), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2093_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2093_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2093_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2093__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_139), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2093__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_139), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2093__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_139), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2093__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_139), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2093__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_139), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2093__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_139), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2093__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module AVG_SPEED_U9
//

module AVG_SPEED_U9 (\speed_avg_m3[0] , clk_1mhz, \speed_m3[0] , \speed_avg_m3[1] , 
            \speed_m3[1] , \speed_avg_m3[2] , \speed_m3[2] , \speed_avg_m3[3] , 
            \speed_m3[3] , \speed_avg_m3[4] , \speed_m3[4] , \speed_avg_m3[5] , 
            \speed_m3[5] , \speed_avg_m3[6] , \speed_m3[6] , \speed_avg_m3[7] , 
            \speed_m3[7] , \speed_avg_m3[8] , \speed_m3[8] , \speed_avg_m3[9] , 
            \speed_m3[9] , \speed_avg_m3[10] , \speed_m3[10] , \speed_avg_m3[11] , 
            \speed_m3[11] , \speed_avg_m3[12] , \speed_m3[12] , \speed_avg_m3[13] , 
            \speed_m3[13] , \speed_avg_m3[14] , \speed_m3[14] , \speed_avg_m3[15] , 
            \speed_m3[15] , \speed_avg_m3[16] , \speed_m3[16] , \speed_avg_m3[17] , 
            \speed_m3[17] , \speed_avg_m3[18] , \speed_m3[18] , \speed_avg_m3[19] , 
            \speed_m3[19] , GND_net);
    output \speed_avg_m3[0] ;
    input clk_1mhz;
    input \speed_m3[0] ;
    output \speed_avg_m3[1] ;
    input \speed_m3[1] ;
    output \speed_avg_m3[2] ;
    input \speed_m3[2] ;
    output \speed_avg_m3[3] ;
    input \speed_m3[3] ;
    output \speed_avg_m3[4] ;
    input \speed_m3[4] ;
    output \speed_avg_m3[5] ;
    input \speed_m3[5] ;
    output \speed_avg_m3[6] ;
    input \speed_m3[6] ;
    output \speed_avg_m3[7] ;
    input \speed_m3[7] ;
    output \speed_avg_m3[8] ;
    input \speed_m3[8] ;
    output \speed_avg_m3[9] ;
    input \speed_m3[9] ;
    output \speed_avg_m3[10] ;
    input \speed_m3[10] ;
    output \speed_avg_m3[11] ;
    input \speed_m3[11] ;
    output \speed_avg_m3[12] ;
    input \speed_m3[12] ;
    output \speed_avg_m3[13] ;
    input \speed_m3[13] ;
    output \speed_avg_m3[14] ;
    input \speed_m3[14] ;
    output \speed_avg_m3[15] ;
    input \speed_m3[15] ;
    output \speed_avg_m3[16] ;
    input \speed_m3[16] ;
    output \speed_avg_m3[17] ;
    input \speed_m3[17] ;
    output \speed_avg_m3[18] ;
    input \speed_m3[18] ;
    output \speed_avg_m3[19] ;
    input \speed_m3[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_120;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n19776, n6, n18188, n18187, n18186;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m3[0] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2091__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_120), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091__i0.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m3[1] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m3[2] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m3[3] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m3[4] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m3[5] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m3[6] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m3[7] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m3[8] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m3[9] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m3[10] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m3[11] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m3[12] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m3[13] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m3[14] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m3[15] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m3[16] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m3[17] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m3[18] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m3[19] ), .SP(clk_1mhz_enable_120), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    LUT4 i17187_4_lut (.A(clk_cnt[0]), .B(n19776), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_120)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17187_4_lut.init = 16'h0004;
    LUT4 i16387_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n19776)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16387_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    CCU2D clk_cnt_2091_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18188), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2091_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2091_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2091_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2091_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18187), .COUT(n18188), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2091_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2091_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2091_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2091_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18186), .COUT(n18187), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2091_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2091_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2091_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2091_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18186), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2091_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2091_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2091_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2091__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_120), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2091__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_120), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2091__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_120), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2091__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_120), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2091__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_120), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2091__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_120), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2091__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module AVG_SPEED_U10
//

module AVG_SPEED_U10 (\speed_avg_m2[0] , clk_1mhz, \speed_m2[0] , \speed_avg_m2[1] , 
            \speed_m2[1] , \speed_avg_m2[2] , \speed_m2[2] , \speed_avg_m2[3] , 
            \speed_m2[3] , \speed_avg_m2[4] , \speed_m2[4] , \speed_avg_m2[5] , 
            \speed_m2[5] , \speed_avg_m2[6] , \speed_m2[6] , \speed_avg_m2[7] , 
            \speed_m2[7] , \speed_avg_m2[8] , \speed_m2[8] , \speed_avg_m2[9] , 
            \speed_m2[9] , \speed_avg_m2[10] , \speed_m2[10] , \speed_avg_m2[11] , 
            \speed_m2[11] , \speed_avg_m2[12] , \speed_m2[12] , \speed_avg_m2[13] , 
            \speed_m2[13] , \speed_avg_m2[14] , \speed_m2[14] , \speed_avg_m2[15] , 
            \speed_m2[15] , \speed_avg_m2[16] , \speed_m2[16] , \speed_avg_m2[17] , 
            \speed_m2[17] , \speed_avg_m2[18] , \speed_m2[18] , \speed_avg_m2[19] , 
            \speed_m2[19] , GND_net);
    output \speed_avg_m2[0] ;
    input clk_1mhz;
    input \speed_m2[0] ;
    output \speed_avg_m2[1] ;
    input \speed_m2[1] ;
    output \speed_avg_m2[2] ;
    input \speed_m2[2] ;
    output \speed_avg_m2[3] ;
    input \speed_m2[3] ;
    output \speed_avg_m2[4] ;
    input \speed_m2[4] ;
    output \speed_avg_m2[5] ;
    input \speed_m2[5] ;
    output \speed_avg_m2[6] ;
    input \speed_m2[6] ;
    output \speed_avg_m2[7] ;
    input \speed_m2[7] ;
    output \speed_avg_m2[8] ;
    input \speed_m2[8] ;
    output \speed_avg_m2[9] ;
    input \speed_m2[9] ;
    output \speed_avg_m2[10] ;
    input \speed_m2[10] ;
    output \speed_avg_m2[11] ;
    input \speed_m2[11] ;
    output \speed_avg_m2[12] ;
    input \speed_m2[12] ;
    output \speed_avg_m2[13] ;
    input \speed_m2[13] ;
    output \speed_avg_m2[14] ;
    input \speed_m2[14] ;
    output \speed_avg_m2[15] ;
    input \speed_m2[15] ;
    output \speed_avg_m2[16] ;
    input \speed_m2[16] ;
    output \speed_avg_m2[17] ;
    input \speed_m2[17] ;
    output \speed_avg_m2[18] ;
    input \speed_m2[18] ;
    output \speed_avg_m2[19] ;
    input \speed_m2[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_101;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n19778, n6, n18192, n18191, n18190;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m2[0] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2089__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_101), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089__i0.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m2[1] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m2[2] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m2[3] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m2[4] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m2[5] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m2[6] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m2[7] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m2[8] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m2[9] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m2[10] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m2[11] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m2[12] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m2[13] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m2[14] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m2[15] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m2[16] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m2[17] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m2[18] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m2[19] ), .SP(clk_1mhz_enable_101), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    LUT4 i17193_4_lut (.A(clk_cnt[0]), .B(n19778), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_101)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17193_4_lut.init = 16'h0004;
    LUT4 i16389_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n19778)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16389_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    CCU2D clk_cnt_2089_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18192), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2089_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2089_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2089_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2089_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18191), .COUT(n18192), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2089_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2089_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2089_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2089_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18190), .COUT(n18191), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2089_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2089_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2089_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2089_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18190), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2089_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2089_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2089_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2089__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_101), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2089__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_101), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2089__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_101), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2089__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_101), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2089__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_101), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2089__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_101), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2089__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AVG_SPEED_U11
//

module AVG_SPEED_U11 (\speed_avg_m1[0] , clk_1mhz, \speed_m1[0] , \speed_avg_m1[1] , 
            \speed_m1[1] , \speed_avg_m1[2] , \speed_m1[2] , \speed_avg_m1[3] , 
            \speed_m1[3] , \speed_avg_m1[4] , \speed_m1[4] , \speed_avg_m1[5] , 
            \speed_m1[5] , \speed_avg_m1[6] , \speed_m1[6] , \speed_avg_m1[7] , 
            \speed_m1[7] , \speed_avg_m1[8] , \speed_m1[8] , \speed_avg_m1[9] , 
            \speed_m1[9] , \speed_avg_m1[10] , \speed_m1[10] , \speed_avg_m1[11] , 
            \speed_m1[11] , \speed_avg_m1[12] , \speed_m1[12] , \speed_avg_m1[13] , 
            \speed_m1[13] , \speed_avg_m1[14] , \speed_m1[14] , \speed_avg_m1[15] , 
            \speed_m1[15] , \speed_avg_m1[16] , \speed_m1[16] , \speed_avg_m1[17] , 
            \speed_m1[17] , \speed_avg_m1[18] , \speed_m1[18] , \speed_avg_m1[19] , 
            \speed_m1[19] , GND_net);
    output \speed_avg_m1[0] ;
    input clk_1mhz;
    input \speed_m1[0] ;
    output \speed_avg_m1[1] ;
    input \speed_m1[1] ;
    output \speed_avg_m1[2] ;
    input \speed_m1[2] ;
    output \speed_avg_m1[3] ;
    input \speed_m1[3] ;
    output \speed_avg_m1[4] ;
    input \speed_m1[4] ;
    output \speed_avg_m1[5] ;
    input \speed_m1[5] ;
    output \speed_avg_m1[6] ;
    input \speed_m1[6] ;
    output \speed_avg_m1[7] ;
    input \speed_m1[7] ;
    output \speed_avg_m1[8] ;
    input \speed_m1[8] ;
    output \speed_avg_m1[9] ;
    input \speed_m1[9] ;
    output \speed_avg_m1[10] ;
    input \speed_m1[10] ;
    output \speed_avg_m1[11] ;
    input \speed_m1[11] ;
    output \speed_avg_m1[12] ;
    input \speed_m1[12] ;
    output \speed_avg_m1[13] ;
    input \speed_m1[13] ;
    output \speed_avg_m1[14] ;
    input \speed_m1[14] ;
    output \speed_avg_m1[15] ;
    input \speed_m1[15] ;
    output \speed_avg_m1[16] ;
    input \speed_m1[16] ;
    output \speed_avg_m1[17] ;
    input \speed_m1[17] ;
    output \speed_avg_m1[18] ;
    input \speed_m1[18] ;
    output \speed_avg_m1[19] ;
    input \speed_m1[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_82;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n12, n18196, n18195, n18194;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m1[0] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2087__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_82), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087__i0.GSR = "DISABLED";
    LUT4 i17190_4_lut (.A(clk_cnt[2]), .B(n12), .C(clk_cnt[1]), .D(clk_cnt[6]), 
         .Z(clk_1mhz_enable_82)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17190_4_lut.init = 16'h0200;
    LUT4 i5_4_lut (.A(clk_cnt[4]), .B(clk_cnt[3]), .C(clk_cnt[0]), .D(clk_cnt[5]), 
         .Z(n12)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i5_4_lut.init = 16'hfeff;
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m1[1] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m1[2] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m1[3] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m1[4] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m1[5] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m1[6] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m1[7] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m1[8] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m1[9] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m1[10] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m1[11] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m1[12] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m1[13] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m1[14] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m1[15] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m1[16] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m1[17] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m1[18] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m1[19] ), .SP(clk_1mhz_enable_82), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    CCU2D clk_cnt_2087_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18196), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2087_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2087_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2087_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2087_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18195), .COUT(n18196), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2087_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2087_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2087_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2087_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18194), .COUT(n18195), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2087_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2087_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2087_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2087_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18194), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2087_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2087_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2087_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2087__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_82), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2087__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_82), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2087__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_82), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2087__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_82), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2087__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_82), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2087__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_82), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2087__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module SPI
//

module SPI (GND_net, speed_set_m4, clkout_c, MISO_N_624, clkout_c_enable_172, 
            enable_m1, enable_m2, enable_m3, enable_m4, clkout_c_enable_173, 
            CS_c, SCK_c, speed_set_m3, hallsense_m1, dir_m1, n2860, 
            n2896, hallsense_m2, dir_m2, n2968, n3004, rst, MOSI_c, 
            hallsense_m3, dir_m3, n3076, n3112, n22100, n21354, 
            hallsense_m4, dir_m4, n3184, n3220, \send_buffer[94] , 
            \send_buffer_95__N_346[94] , \speed_avg_m1[0] , \speed_avg_m1[8] , 
            \speed_avg_m1[9] , \speed_avg_m2[19] , \speed_avg_m1[10] , 
            \speed_avg_m1[6] , \speed_avg_m1[7] , \speed_avg_m1[4] , \speed_avg_m1[2] , 
            \speed_avg_m1[1] , \speed_avg_m1[3] , \speed_avg_m1[5] , \speed_avg_m1[11] , 
            \speed_avg_m1[12] , \speed_avg_m1[13] , \speed_avg_m1[14] , 
            \speed_avg_m1[15] , \speed_avg_m1[16] , \speed_avg_m1[17] , 
            \speed_avg_m1[18] , \speed_avg_m4[8] , \speed_avg_m4[7] , 
            \speed_avg_m4[10] , \speed_avg_m4[9] , \speed_avg_m4[11] , 
            \speed_avg_m4[12] , \speed_avg_m4[13] , \speed_avg_m4[14] , 
            \speed_avg_m4[15] , \speed_avg_m4[16] , \speed_avg_m4[17] , 
            \speed_avg_m4[18] , \speed_avg_m4[19] , \speed_avg_m3[0] , 
            \speed_avg_m3[1] , \speed_avg_m3[2] , \speed_avg_m3[3] , \speed_avg_m3[4] , 
            \speed_avg_m3[5] , \speed_avg_m3[6] , \speed_avg_m3[7] , \speed_avg_m3[8] , 
            \speed_avg_m3[9] , \speed_avg_m3[10] , \speed_avg_m3[11] , 
            speed_set_m2, \speed_avg_m3[12] , \speed_avg_m3[13] , \speed_avg_m3[14] , 
            speed_set_m1, \speed_avg_m3[15] , \speed_avg_m3[16] , \speed_avg_m3[17] , 
            \speed_avg_m3[18] , \speed_avg_m3[19] , \speed_avg_m2[0] , 
            \speed_avg_m2[1] , \speed_avg_m2[2] , \speed_avg_m2[3] , \speed_avg_m2[4] , 
            \speed_avg_m2[5] , \speed_avg_m2[6] , \speed_avg_m2[7] , \speed_avg_m2[8] , 
            \speed_avg_m2[9] , \speed_avg_m2[10] , \speed_avg_m2[11] , 
            \speed_avg_m2[12] , \speed_avg_m2[13] , \speed_avg_m2[14] , 
            \speed_avg_m2[15] , \speed_avg_m2[16] , \speed_avg_m2[17] , 
            \speed_avg_m2[18] , \speed_avg_m4[0] , \speed_avg_m4[1] , 
            \speed_avg_m1[19] , \speed_avg_m4[2] , \speed_avg_m4[3] , 
            \speed_avg_m4[4] , \speed_avg_m4[5] , \speed_avg_m4[6] , n21336, 
            n5132, free_m4, n19415, free_m3, n19427, free_m2, n19411, 
            free_m1, n19421);
    input GND_net;
    output [20:0]speed_set_m4;
    input clkout_c;
    output MISO_N_624;
    input clkout_c_enable_172;
    output enable_m1;
    output enable_m2;
    output enable_m3;
    output enable_m4;
    input clkout_c_enable_173;
    input CS_c;
    input SCK_c;
    output [20:0]speed_set_m3;
    input [2:0]hallsense_m1;
    input dir_m1;
    output n2860;
    output n2896;
    input [2:0]hallsense_m2;
    input dir_m2;
    output n2968;
    output n3004;
    input rst;
    input MOSI_c;
    input [2:0]hallsense_m3;
    input dir_m3;
    output n3076;
    output n3112;
    input n22100;
    output n21354;
    input [2:0]hallsense_m4;
    input dir_m4;
    output n3184;
    output n3220;
    output \send_buffer[94] ;
    input \send_buffer_95__N_346[94] ;
    input \speed_avg_m1[0] ;
    input \speed_avg_m1[8] ;
    input \speed_avg_m1[9] ;
    input \speed_avg_m2[19] ;
    input \speed_avg_m1[10] ;
    input \speed_avg_m1[6] ;
    input \speed_avg_m1[7] ;
    input \speed_avg_m1[4] ;
    input \speed_avg_m1[2] ;
    input \speed_avg_m1[1] ;
    input \speed_avg_m1[3] ;
    input \speed_avg_m1[5] ;
    input \speed_avg_m1[11] ;
    input \speed_avg_m1[12] ;
    input \speed_avg_m1[13] ;
    input \speed_avg_m1[14] ;
    input \speed_avg_m1[15] ;
    input \speed_avg_m1[16] ;
    input \speed_avg_m1[17] ;
    input \speed_avg_m1[18] ;
    input \speed_avg_m4[8] ;
    input \speed_avg_m4[7] ;
    input \speed_avg_m4[10] ;
    input \speed_avg_m4[9] ;
    input \speed_avg_m4[11] ;
    input \speed_avg_m4[12] ;
    input \speed_avg_m4[13] ;
    input \speed_avg_m4[14] ;
    input \speed_avg_m4[15] ;
    input \speed_avg_m4[16] ;
    input \speed_avg_m4[17] ;
    input \speed_avg_m4[18] ;
    input \speed_avg_m4[19] ;
    input \speed_avg_m3[0] ;
    input \speed_avg_m3[1] ;
    input \speed_avg_m3[2] ;
    input \speed_avg_m3[3] ;
    input \speed_avg_m3[4] ;
    input \speed_avg_m3[5] ;
    input \speed_avg_m3[6] ;
    input \speed_avg_m3[7] ;
    input \speed_avg_m3[8] ;
    input \speed_avg_m3[9] ;
    input \speed_avg_m3[10] ;
    input \speed_avg_m3[11] ;
    output [20:0]speed_set_m2;
    input \speed_avg_m3[12] ;
    input \speed_avg_m3[13] ;
    input \speed_avg_m3[14] ;
    output [20:0]speed_set_m1;
    input \speed_avg_m3[15] ;
    input \speed_avg_m3[16] ;
    input \speed_avg_m3[17] ;
    input \speed_avg_m3[18] ;
    input \speed_avg_m3[19] ;
    input \speed_avg_m2[0] ;
    input \speed_avg_m2[1] ;
    input \speed_avg_m2[2] ;
    input \speed_avg_m2[3] ;
    input \speed_avg_m2[4] ;
    input \speed_avg_m2[5] ;
    input \speed_avg_m2[6] ;
    input \speed_avg_m2[7] ;
    input \speed_avg_m2[8] ;
    input \speed_avg_m2[9] ;
    input \speed_avg_m2[10] ;
    input \speed_avg_m2[11] ;
    input \speed_avg_m2[12] ;
    input \speed_avg_m2[13] ;
    input \speed_avg_m2[14] ;
    input \speed_avg_m2[15] ;
    input \speed_avg_m2[16] ;
    input \speed_avg_m2[17] ;
    input \speed_avg_m2[18] ;
    input \speed_avg_m4[0] ;
    input \speed_avg_m4[1] ;
    input \speed_avg_m1[19] ;
    input \speed_avg_m4[2] ;
    input \speed_avg_m4[3] ;
    input \speed_avg_m4[4] ;
    input \speed_avg_m4[5] ;
    input \speed_avg_m4[6] ;
    output n21336;
    output n5132;
    input free_m4;
    output n19415;
    input free_m3;
    output n19427;
    input free_m2;
    output n19411;
    input free_m1;
    output n19421;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire n18288;
    wire [95:0]recv_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(68[10:21])
    
    wire n18289, clkout_c_enable_254, n14142, MISO_N_670, n18287, 
        n18286, n18285, n18284, n18283, n18282, n18281, n18280, 
        n18279, n3388, n18278, n18277, MISOb, MISOb_N_660, enable_m1_N_633, 
        enable_m1_N_627;
    wire [83:0]n169;
    
    wire enable_m2_N_635, enable_m3_N_642, enable_m4_N_649, CSold, CSlatched, 
        SCKold, SCKlatched;
    wire [95:0]send_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(67[10:21])
    
    wire n21386, n18276, n18275, n18274, n14162, n18273, n21385, 
        MISO_N_625, CSlatched_N_664, n18272, n21374, clkout_c_enable_60, 
        n22086, n22087, n21355;
    wire [95:0]send_buffer_95__N_346;
    
    wire n21370, n22098;
    wire [95:0]MISOb_N_666;
    
    wire n21289, n22090, n22091, clkout_c_enable_94, n21365, n21288, 
        n21360, n21335, n3340, n3316, n39_adj_2202, n40_adj_2203, 
        n36_adj_2204, n28_adj_2205, n38_adj_2206, n32_adj_2207, n34_adj_2208, 
        n24_adj_2209, n3364, n39_adj_2210, n40_adj_2211, n36_adj_2212, 
        n28_adj_2213, n38_adj_2214, n32_adj_2215, n34_adj_2216, n24_adj_2217, 
        n3436, n3412, n39_adj_2218, n40_adj_2219, n36_adj_2220, n28_adj_2221, 
        n38_adj_2222, n32_adj_2223, n3484, n3460, n39_adj_2224, n40_adj_2225, 
        n34_adj_2226, n24_adj_2227, n36_adj_2228, n28_adj_2229, n38_adj_2230, 
        n32_adj_2231, n18271, n18270, n14202, n14182, n18269, n18268, 
        n18267, n34_adj_2232, n24_adj_2233, n18266, n18265, n18264, 
        n18263, n18262, n18261, n18260, n18259, n18102, n18258, 
        n18101, n18100, n18257, n18099, n18256, n18255, n18254, 
        n18098, n18097, n18096, n18095, n18094, n18093, n18307, 
        n18306, n18072, n18305, n18304, n18071, n18070, n18069, 
        n18068, n18303, n18302, n18301, n18300, n18067, n18299, 
        n18066, n18298, n18297, n18296, n18065, n18295, n18294, 
        n18293, n18292, n18291, n18290;
    
    CCU2D add_15009_19 (.A0(recv_buffer[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18288), .COUT(n18289));
    defparam add_15009_19.INIT0 = 16'hf555;
    defparam add_15009_19.INIT1 = 16'hf555;
    defparam add_15009_19.INJECT1_0 = "NO";
    defparam add_15009_19.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i20 (.D(recv_buffer[32]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i20.GSR = "DISABLED";
    FD1S3AX MISO_124 (.D(MISO_N_670), .CK(clkout_c), .Q(MISO_N_624)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISO_124.GSR = "DISABLED";
    CCU2D add_15009_17 (.A0(recv_buffer[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18287), .COUT(n18288));
    defparam add_15009_17.INIT0 = 16'hf555;
    defparam add_15009_17.INIT1 = 16'hf555;
    defparam add_15009_17.INJECT1_0 = "NO";
    defparam add_15009_17.INJECT1_1 = "NO";
    CCU2D add_15009_15 (.A0(recv_buffer[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18286), .COUT(n18287));
    defparam add_15009_15.INIT0 = 16'hf555;
    defparam add_15009_15.INIT1 = 16'hf555;
    defparam add_15009_15.INJECT1_0 = "NO";
    defparam add_15009_15.INJECT1_1 = "NO";
    CCU2D add_15009_13 (.A0(recv_buffer[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18285), .COUT(n18286));
    defparam add_15009_13.INIT0 = 16'hf555;
    defparam add_15009_13.INIT1 = 16'h0aaa;
    defparam add_15009_13.INJECT1_0 = "NO";
    defparam add_15009_13.INJECT1_1 = "NO";
    CCU2D add_15009_11 (.A0(recv_buffer[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18284), .COUT(n18285));
    defparam add_15009_11.INIT0 = 16'h0aaa;
    defparam add_15009_11.INIT1 = 16'hf555;
    defparam add_15009_11.INJECT1_0 = "NO";
    defparam add_15009_11.INJECT1_1 = "NO";
    CCU2D add_15009_9 (.A0(recv_buffer[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18283), .COUT(n18284));
    defparam add_15009_9.INIT0 = 16'h0aaa;
    defparam add_15009_9.INIT1 = 16'h0aaa;
    defparam add_15009_9.INJECT1_0 = "NO";
    defparam add_15009_9.INJECT1_1 = "NO";
    CCU2D add_15009_7 (.A0(recv_buffer[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18282), .COUT(n18283));
    defparam add_15009_7.INIT0 = 16'hf555;
    defparam add_15009_7.INIT1 = 16'hf555;
    defparam add_15009_7.INJECT1_0 = "NO";
    defparam add_15009_7.INJECT1_1 = "NO";
    CCU2D add_15009_5 (.A0(recv_buffer[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18281), .COUT(n18282));
    defparam add_15009_5.INIT0 = 16'h0aaa;
    defparam add_15009_5.INIT1 = 16'hf555;
    defparam add_15009_5.INJECT1_0 = "NO";
    defparam add_15009_5.INJECT1_1 = "NO";
    CCU2D add_15009_3 (.A0(recv_buffer[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18280), .COUT(n18281));
    defparam add_15009_3.INIT0 = 16'hf555;
    defparam add_15009_3.INIT1 = 16'hf555;
    defparam add_15009_3.INJECT1_0 = "NO";
    defparam add_15009_3.INJECT1_1 = "NO";
    CCU2D add_15009_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[33]), .B1(recv_buffer[34]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18280));
    defparam add_15009_1.INIT0 = 16'hF000;
    defparam add_15009_1.INIT1 = 16'ha666;
    defparam add_15009_1.INJECT1_0 = "NO";
    defparam add_15009_1.INJECT1_1 = "NO";
    CCU2D add_15010_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18279), 
          .S0(n3388));
    defparam add_15010_cout.INIT0 = 16'h0000;
    defparam add_15010_cout.INIT1 = 16'h0000;
    defparam add_15010_cout.INJECT1_0 = "NO";
    defparam add_15010_cout.INJECT1_1 = "NO";
    CCU2D add_15010_16 (.A0(recv_buffer[73]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[74]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18278), .COUT(n18279));
    defparam add_15010_16.INIT0 = 16'h5aaa;
    defparam add_15010_16.INIT1 = 16'h0aaa;
    defparam add_15010_16.INJECT1_0 = "NO";
    defparam add_15010_16.INJECT1_1 = "NO";
    CCU2D add_15010_14 (.A0(recv_buffer[71]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[72]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18277), .COUT(n18278));
    defparam add_15010_14.INIT0 = 16'h5aaa;
    defparam add_15010_14.INIT1 = 16'h5aaa;
    defparam add_15010_14.INJECT1_0 = "NO";
    defparam add_15010_14.INJECT1_1 = "NO";
    FD1P3AX MISOb_118 (.D(MISOb_N_660), .SP(clkout_c_enable_172), .CK(clkout_c), 
            .Q(MISOb));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISOb_118.GSR = "DISABLED";
    FD1P3AX enable_m1_109 (.D(enable_m1_N_627), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m1_109.GSR = "ENABLED";
    FD1P3IX speed_set_m4_i0_i0 (.D(n169[0]), .SP(clkout_c_enable_254), .CD(n14142), 
            .CK(clkout_c), .Q(speed_set_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i0.GSR = "DISABLED";
    FD1P3AX enable_m2_110 (.D(enable_m2_N_635), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m2_110.GSR = "ENABLED";
    FD1P3AX enable_m3_111 (.D(enable_m3_N_642), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m3_111.GSR = "ENABLED";
    FD1P3AX enable_m4_112 (.D(enable_m4_N_649), .SP(enable_m1_N_633), .CK(clkout_c), 
            .Q(enable_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m4_112.GSR = "ENABLED";
    FD1P3AX CSold_113 (.D(CSlatched), .SP(clkout_c_enable_173), .CK(clkout_c), 
            .Q(CSold));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_113.GSR = "DISABLED";
    FD1P3AX SCKold_114 (.D(SCKlatched), .SP(clkout_c_enable_173), .CK(clkout_c), 
            .Q(SCKold));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKold_114.GSR = "DISABLED";
    FD1P3AX CSlatched_115 (.D(CS_c), .SP(clkout_c_enable_173), .CK(clkout_c), 
            .Q(CSlatched));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_115.GSR = "DISABLED";
    FD1P3AX SCKlatched_116 (.D(SCK_c), .SP(clkout_c_enable_173), .CK(clkout_c), 
            .Q(SCKlatched));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKlatched_116.GSR = "DISABLED";
    LUT4 i2933_3_lut_4_lut_then_4_lut (.A(CSlatched), .B(MISOb), .C(CSold), 
         .D(send_buffer[1]), .Z(n21386)) /* synthesis lut_function=(A (B)+!A (C+(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam i2933_3_lut_4_lut_then_4_lut.init = 16'hddd8;
    CCU2D add_15010_12 (.A0(recv_buffer[69]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[70]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18276), .COUT(n18277));
    defparam add_15010_12.INIT0 = 16'h5aaa;
    defparam add_15010_12.INIT1 = 16'h5aaa;
    defparam add_15010_12.INJECT1_0 = "NO";
    defparam add_15010_12.INJECT1_1 = "NO";
    CCU2D add_15010_10 (.A0(recv_buffer[67]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[68]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18275), .COUT(n18276));
    defparam add_15010_10.INIT0 = 16'h5555;
    defparam add_15010_10.INIT1 = 16'h5aaa;
    defparam add_15010_10.INJECT1_0 = "NO";
    defparam add_15010_10.INJECT1_1 = "NO";
    CCU2D add_15010_8 (.A0(recv_buffer[65]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[66]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18274), .COUT(n18275));
    defparam add_15010_8.INIT0 = 16'h5aaa;
    defparam add_15010_8.INIT1 = 16'h5aaa;
    defparam add_15010_8.INJECT1_0 = "NO";
    defparam add_15010_8.INJECT1_1 = "NO";
    FD1P3IX speed_set_m3_i0_i0 (.D(recv_buffer[33]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i0.GSR = "DISABLED";
    CCU2D add_15010_6 (.A0(recv_buffer[63]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[64]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18273), .COUT(n18274));
    defparam add_15010_6.INIT0 = 16'h5555;
    defparam add_15010_6.INIT1 = 16'h5555;
    defparam add_15010_6.INJECT1_0 = "NO";
    defparam add_15010_6.INJECT1_1 = "NO";
    LUT4 i2933_3_lut_4_lut_else_4_lut (.A(CSlatched), .B(MISOb), .C(CSold), 
         .Z(n21385)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam i2933_3_lut_4_lut_else_4_lut.init = 16'h8c8c;
    FD1P3AX i101_125 (.D(CSlatched_N_664), .SP(clkout_c_enable_173), .CK(clkout_c), 
            .Q(MISO_N_625));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i101_125.GSR = "DISABLED";
    CCU2D add_15010_4 (.A0(recv_buffer[61]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[62]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18272), .COUT(n18273));
    defparam add_15010_4.INIT0 = 16'h5aaa;
    defparam add_15010_4.INIT1 = 16'h5555;
    defparam add_15010_4.INJECT1_0 = "NO";
    defparam add_15010_4.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(hallsense_m1[2]), .B(n21374), .C(dir_m1), .D(hallsense_m1[1]), 
         .Z(n2860)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut.init = 16'h4008;
    LUT4 i1_4_lut_adj_133 (.A(hallsense_m1[1]), .B(n21374), .C(dir_m1), 
         .D(hallsense_m1[0]), .Z(n2896)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_133.init = 16'h4008;
    FD1P3AX \SPI__5_rep_5__i0  (.D(recv_buffer[13]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(n169[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5_rep_5__i0 .GSR = "DISABLED";
    PFUMX i17483 (.BLUT(n22086), .ALUT(n22087), .C0(n21355), .Z(send_buffer_95__N_346[1]));
    LUT4 i1_4_lut_adj_134 (.A(hallsense_m2[2]), .B(n21370), .C(dir_m2), 
         .D(hallsense_m2[1]), .Z(n2968)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_134.init = 16'h4008;
    LUT4 i1_4_lut_adj_135 (.A(hallsense_m2[1]), .B(n21370), .C(dir_m2), 
         .D(hallsense_m2[0]), .Z(n3004)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_135.init = 16'h4008;
    PFUMX i17313 (.BLUT(n21385), .ALUT(n21386), .C0(n21355), .Z(MISOb_N_660));
    FD1P3AX CSold_113_rep_407 (.D(CSlatched), .SP(rst), .CK(clkout_c), 
            .Q(n22098));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_113_rep_407.GSR = "DISABLED";
    LUT4 mux_51_i5_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[5]), 
         .D(MISOb_N_666[4]), .Z(send_buffer_95__N_346[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i7_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[7]), 
         .D(MISOb_N_666[6]), .Z(send_buffer_95__N_346[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i6_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[6]), 
         .D(MISOb_N_666[5]), .Z(send_buffer_95__N_346[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i8_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[8]), 
         .D(MISOb_N_666[7]), .Z(send_buffer_95__N_346[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i9_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[9]), 
         .D(MISOb_N_666[8]), .Z(send_buffer_95__N_346[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i10_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[10]), 
         .D(MISOb_N_666[9]), .Z(send_buffer_95__N_346[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i11_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[11]), 
         .D(MISOb_N_666[10]), .Z(send_buffer_95__N_346[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i12_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[12]), 
         .D(MISOb_N_666[11]), .Z(send_buffer_95__N_346[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i13_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[13]), 
         .D(MISOb_N_666[12]), .Z(send_buffer_95__N_346[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i14_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[14]), 
         .D(MISOb_N_666[13]), .Z(send_buffer_95__N_346[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i15_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[15]), 
         .D(MISOb_N_666[14]), .Z(send_buffer_95__N_346[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i16_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[16]), 
         .D(MISOb_N_666[15]), .Z(send_buffer_95__N_346[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i17_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[17]), 
         .D(MISOb_N_666[16]), .Z(send_buffer_95__N_346[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i18_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[18]), 
         .D(MISOb_N_666[17]), .Z(send_buffer_95__N_346[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 MISOb_N_667_bdd_2_lut (.A(MISO_N_624), .B(MISO_N_625), .Z(n21289)) /* synthesis lut_function=(A (B)) */ ;
    defparam MISOb_N_667_bdd_2_lut.init = 16'h8888;
    LUT4 mux_51_i19_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[19]), 
         .D(MISOb_N_666[18]), .Z(send_buffer_95__N_346[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i20_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[20]), 
         .D(MISOb_N_666[19]), .Z(send_buffer_95__N_346[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i21_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[21]), 
         .D(MISOb_N_666[20]), .Z(send_buffer_95__N_346[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i22_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[22]), 
         .D(MISOb_N_666[21]), .Z(send_buffer_95__N_346[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i23_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[23]), 
         .D(MISOb_N_666[22]), .Z(send_buffer_95__N_346[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i24_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[24]), 
         .D(MISOb_N_666[23]), .Z(send_buffer_95__N_346[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i25_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[25]), 
         .D(MISOb_N_666[24]), .Z(send_buffer_95__N_346[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i25_3_lut_4_lut.init = 16'hfd20;
    PFUMX i17486 (.BLUT(n22090), .ALUT(n22091), .C0(n21355), .Z(send_buffer_95__N_346[2]));
    LUT4 mux_51_i26_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[26]), 
         .D(MISOb_N_666[25]), .Z(send_buffer_95__N_346[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i27_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[27]), 
         .D(MISOb_N_666[26]), .Z(send_buffer_95__N_346[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i28_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[28]), 
         .D(MISOb_N_666[27]), .Z(send_buffer_95__N_346[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i29_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[29]), 
         .D(MISOb_N_666[28]), .Z(send_buffer_95__N_346[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i29_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX \SPI__5__i83  (.D(MOSI_c), .SP(clkout_c_enable_60), .CK(clkout_c), 
            .Q(recv_buffer[95]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i83 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i82  (.D(recv_buffer[95]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[94]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i82 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i81  (.D(recv_buffer[94]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[93]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i81 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i80  (.D(recv_buffer[93]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[92]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i80 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i79  (.D(recv_buffer[92]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[91]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i79 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i78  (.D(recv_buffer[91]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[90]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i78 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i77  (.D(recv_buffer[90]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[89]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i77 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i76  (.D(recv_buffer[89]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[88]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i76 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i75  (.D(recv_buffer[88]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[87]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i75 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i74  (.D(recv_buffer[87]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[86]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i74 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i73  (.D(recv_buffer[86]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[85]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i73 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i72  (.D(recv_buffer[85]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[84]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i72 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i71  (.D(recv_buffer[84]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[83]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i71 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i70  (.D(recv_buffer[83]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[82]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i70 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i69  (.D(recv_buffer[82]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[81]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i69 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i68  (.D(recv_buffer[81]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[80]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i68 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i67  (.D(recv_buffer[80]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[79]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i67 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i66  (.D(recv_buffer[79]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[78]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i66 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i65  (.D(recv_buffer[78]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[77]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i65 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i64  (.D(recv_buffer[77]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[76]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i64 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i63  (.D(recv_buffer[76]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[75]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i63 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i62  (.D(recv_buffer[75]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[74]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i62 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i61  (.D(recv_buffer[74]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[73]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i61 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i60  (.D(recv_buffer[73]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[72]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i60 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i59  (.D(recv_buffer[72]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[71]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i59 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i58  (.D(recv_buffer[71]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[70]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i58 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i57  (.D(recv_buffer[70]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[69]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i57 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i56  (.D(recv_buffer[69]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[68]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i56 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i55  (.D(recv_buffer[68]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[67]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i55 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i54  (.D(recv_buffer[67]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[66]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i54 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i53  (.D(recv_buffer[66]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[65]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i53 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i52  (.D(recv_buffer[65]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[64]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i52 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i51  (.D(recv_buffer[64]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[63]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i51 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i50  (.D(recv_buffer[63]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[62]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i50 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i49  (.D(recv_buffer[62]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[61]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i49 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i48  (.D(recv_buffer[61]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[60]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i48 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i47  (.D(recv_buffer[60]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[59]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i47 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i46  (.D(recv_buffer[59]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[58]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i46 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i45  (.D(recv_buffer[58]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[57]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i45 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i44  (.D(recv_buffer[57]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[56]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i44 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i43  (.D(recv_buffer[56]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[55]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i43 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i42  (.D(recv_buffer[55]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[54]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i42 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i41  (.D(recv_buffer[54]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[53]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i41 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i40  (.D(recv_buffer[53]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[52]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i40 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i39  (.D(recv_buffer[52]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[51]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i39 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i38  (.D(recv_buffer[51]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[50]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i38 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i37  (.D(recv_buffer[50]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[49]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i37 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i36  (.D(recv_buffer[49]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[48]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i36 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i35  (.D(recv_buffer[48]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[47]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i35 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i34  (.D(recv_buffer[47]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[46]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i34 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i33  (.D(recv_buffer[46]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[45]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i33 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i32  (.D(recv_buffer[45]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[44]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i32 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i31  (.D(recv_buffer[44]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[43]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i31 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i30  (.D(recv_buffer[43]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[42]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i30 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i29  (.D(recv_buffer[42]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[41]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i29 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i28  (.D(recv_buffer[41]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[40]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i28 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i27  (.D(recv_buffer[40]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[39]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i27 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i26  (.D(recv_buffer[39]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[38]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i26 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i25  (.D(recv_buffer[38]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[37]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i25 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i24  (.D(recv_buffer[37]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[36]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i24 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i23  (.D(recv_buffer[36]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[35]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i23 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i22  (.D(recv_buffer[35]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[34]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i22 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i21  (.D(recv_buffer[34]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[33]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i21 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i20  (.D(recv_buffer[33]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[32]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i20 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i19  (.D(recv_buffer[32]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[31]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i19 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i18  (.D(recv_buffer[31]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[30]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i18 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i17  (.D(recv_buffer[30]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[29]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i17 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i16  (.D(recv_buffer[29]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[28]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i16 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i15  (.D(recv_buffer[28]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[27]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i15 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i14  (.D(recv_buffer[27]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[26]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i14 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i13  (.D(recv_buffer[26]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[25]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i13 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i12  (.D(recv_buffer[25]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[24]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i12 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i11  (.D(recv_buffer[24]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[23]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i11 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i10  (.D(recv_buffer[23]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[22]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i10 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i9  (.D(recv_buffer[22]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[21]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i9 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i8  (.D(recv_buffer[21]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[20]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i8 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i7  (.D(recv_buffer[20]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i7 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i6  (.D(recv_buffer[19]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i6 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i5  (.D(recv_buffer[18]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[17]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i5 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i4  (.D(recv_buffer[17]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i4 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i3  (.D(recv_buffer[16]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i3 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i2  (.D(recv_buffer[15]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i2 .GSR = "DISABLED";
    FD1P3AX \SPI__5__i1  (.D(recv_buffer[14]), .SP(clkout_c_enable_94), 
            .CK(clkout_c), .Q(recv_buffer[13]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam \SPI__5__i1 .GSR = "DISABLED";
    LUT4 mux_51_i30_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[30]), 
         .D(MISOb_N_666[29]), .Z(send_buffer_95__N_346[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i31_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[31]), 
         .D(MISOb_N_666[30]), .Z(send_buffer_95__N_346[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i31_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i32_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[32]), 
         .D(MISOb_N_666[31]), .Z(send_buffer_95__N_346[31])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i32_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i33_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[33]), 
         .D(MISOb_N_666[32]), .Z(send_buffer_95__N_346[32])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i33_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i34_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[34]), 
         .D(MISOb_N_666[33]), .Z(send_buffer_95__N_346[33])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i34_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i35_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[35]), 
         .D(MISOb_N_666[34]), .Z(send_buffer_95__N_346[34])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i35_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_136 (.A(hallsense_m3[2]), .B(n21365), .C(dir_m3), 
         .D(hallsense_m3[1]), .Z(n3076)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_136.init = 16'h4008;
    LUT4 mux_51_i36_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[36]), 
         .D(MISOb_N_666[35]), .Z(send_buffer_95__N_346[35])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i36_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i37_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[37]), 
         .D(MISOb_N_666[36]), .Z(send_buffer_95__N_346[36])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i37_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i38_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[38]), 
         .D(MISOb_N_666[37]), .Z(send_buffer_95__N_346[37])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i38_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i39_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[39]), 
         .D(MISOb_N_666[38]), .Z(send_buffer_95__N_346[38])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i39_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_137 (.A(hallsense_m3[1]), .B(n21365), .C(dir_m3), 
         .D(hallsense_m3[0]), .Z(n3112)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_137.init = 16'h4008;
    LUT4 mux_51_i40_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[40]), 
         .D(MISOb_N_666[39]), .Z(send_buffer_95__N_346[39])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i40_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i41_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[41]), 
         .D(MISOb_N_666[40]), .Z(send_buffer_95__N_346[40])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i41_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i42_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[42]), 
         .D(MISOb_N_666[41]), .Z(send_buffer_95__N_346[41])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i42_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i43_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[43]), 
         .D(MISOb_N_666[42]), .Z(send_buffer_95__N_346[42])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i43_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i44_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[44]), 
         .D(MISOb_N_666[43]), .Z(send_buffer_95__N_346[43])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i44_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i45_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[45]), 
         .D(MISOb_N_666[44]), .Z(send_buffer_95__N_346[44])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i45_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i46_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[46]), 
         .D(MISOb_N_666[45]), .Z(send_buffer_95__N_346[45])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i46_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i47_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[47]), 
         .D(MISOb_N_666[46]), .Z(send_buffer_95__N_346[46])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i47_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i48_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[48]), 
         .D(MISOb_N_666[47]), .Z(send_buffer_95__N_346[47])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i48_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i49_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[49]), 
         .D(MISOb_N_666[48]), .Z(send_buffer_95__N_346[48])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i49_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i50_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[50]), 
         .D(MISOb_N_666[49]), .Z(send_buffer_95__N_346[49])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i50_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i51_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[51]), 
         .D(MISOb_N_666[50]), .Z(send_buffer_95__N_346[50])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i51_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i52_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[52]), 
         .D(MISOb_N_666[51]), .Z(send_buffer_95__N_346[51])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i52_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i53_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[53]), 
         .D(MISOb_N_666[52]), .Z(send_buffer_95__N_346[52])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i53_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i54_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[54]), 
         .D(MISOb_N_666[53]), .Z(send_buffer_95__N_346[53])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i54_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i55_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[55]), 
         .D(MISOb_N_666[54]), .Z(send_buffer_95__N_346[54])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i55_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i56_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[56]), 
         .D(MISOb_N_666[55]), .Z(send_buffer_95__N_346[55])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i56_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i57_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[57]), 
         .D(MISOb_N_666[56]), .Z(send_buffer_95__N_346[56])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i57_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i58_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[58]), 
         .D(MISOb_N_666[57]), .Z(send_buffer_95__N_346[57])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i58_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i59_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[59]), 
         .D(MISOb_N_666[58]), .Z(send_buffer_95__N_346[58])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i59_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i60_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[60]), 
         .D(MISOb_N_666[59]), .Z(send_buffer_95__N_346[59])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i60_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i61_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[61]), 
         .D(MISOb_N_666[60]), .Z(send_buffer_95__N_346[60])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i61_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i62_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[62]), 
         .D(MISOb_N_666[61]), .Z(send_buffer_95__N_346[61])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i62_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i63_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[63]), 
         .D(MISOb_N_666[62]), .Z(send_buffer_95__N_346[62])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i63_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i64_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[64]), 
         .D(MISOb_N_666[63]), .Z(send_buffer_95__N_346[63])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i64_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3_4_lut_rep_413 (.A(SCKold), .B(n22100), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_60)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut_rep_413.init = 16'h0400;
    LUT4 mux_51_i65_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[65]), 
         .D(MISOb_N_666[64]), .Z(send_buffer_95__N_346[64])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i65_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i66_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[66]), 
         .D(MISOb_N_666[65]), .Z(send_buffer_95__N_346[65])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i66_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i67_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[67]), 
         .D(MISOb_N_666[66]), .Z(send_buffer_95__N_346[66])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i67_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i68_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[68]), 
         .D(MISOb_N_666[67]), .Z(send_buffer_95__N_346[67])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i68_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i69_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[69]), 
         .D(MISOb_N_666[68]), .Z(send_buffer_95__N_346[68])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i69_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i70_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[70]), 
         .D(MISOb_N_666[69]), .Z(send_buffer_95__N_346[69])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i70_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i71_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[71]), 
         .D(MISOb_N_666[70]), .Z(send_buffer_95__N_346[70])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i71_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i72_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[72]), 
         .D(MISOb_N_666[71]), .Z(send_buffer_95__N_346[71])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i72_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i73_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[73]), 
         .D(MISOb_N_666[72]), .Z(send_buffer_95__N_346[72])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i73_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i74_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[74]), 
         .D(MISOb_N_666[73]), .Z(send_buffer_95__N_346[73])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i74_3_lut_4_lut.init = 16'hfd20;
    LUT4 MISOb_N_667_bdd_4_lut (.A(n21355), .B(send_buffer[1]), .C(MISOb), 
         .D(n21354), .Z(n21288)) /* synthesis lut_function=(A (B+(D))+!A !((D)+!C)) */ ;
    defparam MISOb_N_667_bdd_4_lut.init = 16'haad8;
    LUT4 mux_51_i75_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[75]), 
         .D(MISOb_N_666[74]), .Z(send_buffer_95__N_346[74])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i75_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i76_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[76]), 
         .D(MISOb_N_666[75]), .Z(send_buffer_95__N_346[75])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i76_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i77_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[77]), 
         .D(MISOb_N_666[76]), .Z(send_buffer_95__N_346[76])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i77_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i78_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[78]), 
         .D(MISOb_N_666[77]), .Z(send_buffer_95__N_346[77])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i78_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i79_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[79]), 
         .D(MISOb_N_666[78]), .Z(send_buffer_95__N_346[78])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i79_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i80_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[80]), 
         .D(MISOb_N_666[79]), .Z(send_buffer_95__N_346[79])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i80_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_138 (.A(hallsense_m4[2]), .B(n21360), .C(dir_m4), 
         .D(hallsense_m4[1]), .Z(n3184)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_138.init = 16'h4008;
    LUT4 mux_51_i81_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[81]), 
         .D(MISOb_N_666[80]), .Z(send_buffer_95__N_346[80])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i81_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i82_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[82]), 
         .D(MISOb_N_666[81]), .Z(send_buffer_95__N_346[81])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i82_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i83_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[83]), 
         .D(MISOb_N_666[82]), .Z(send_buffer_95__N_346[82])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i83_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i84_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[84]), 
         .D(MISOb_N_666[83]), .Z(send_buffer_95__N_346[83])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i84_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i85_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[85]), 
         .D(MISOb_N_666[84]), .Z(send_buffer_95__N_346[84])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i85_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_139 (.A(hallsense_m4[1]), .B(n21360), .C(dir_m4), 
         .D(hallsense_m4[0]), .Z(n3220)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_4_lut_adj_139.init = 16'h4008;
    LUT4 mux_51_i86_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[86]), 
         .D(MISOb_N_666[85]), .Z(send_buffer_95__N_346[85])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i86_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i87_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[87]), 
         .D(MISOb_N_666[86]), .Z(send_buffer_95__N_346[86])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i87_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i88_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[88]), 
         .D(MISOb_N_666[87]), .Z(send_buffer_95__N_346[87])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i88_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i89_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[89]), 
         .D(MISOb_N_666[88]), .Z(send_buffer_95__N_346[88])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i89_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i90_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[90]), 
         .D(MISOb_N_666[89]), .Z(send_buffer_95__N_346[89])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i90_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i91_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[91]), 
         .D(MISOb_N_666[90]), .Z(send_buffer_95__N_346[90])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i91_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i92_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[92]), 
         .D(MISOb_N_666[91]), .Z(send_buffer_95__N_346[91])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i92_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i93_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[93]), 
         .D(MISOb_N_666[92]), .Z(send_buffer_95__N_346[92])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i93_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i94_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(n21335), 
         .D(MISOb_N_666[93]), .Z(send_buffer_95__N_346[93])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i94_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i4_3_lut_4_lut (.A(n21355), .B(CSlatched), .C(MISOb_N_666[4]), 
         .D(MISOb_N_666[3]), .Z(send_buffer_95__N_346[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_51_i2_3_lut_4_lut_then_4_lut (.A(CSlatched), .B(send_buffer[1]), 
         .C(CSold), .D(send_buffer[2]), .Z(n22087)) /* synthesis lut_function=(A (B)+!A !(C+!(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i2_3_lut_4_lut_then_4_lut.init = 16'h8d88;
    LUT4 CSold_I_0_132_2_lut (.A(CSold), .B(CSlatched), .Z(enable_m1_N_633)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam CSold_I_0_132_2_lut.init = 16'h8888;
    LUT4 i2_4_lut (.A(n3340), .B(n3316), .C(n39_adj_2202), .D(n40_adj_2203), 
         .Z(enable_m1_N_627)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i18_4_lut (.A(recv_buffer[88]), .B(n36_adj_2204), .C(n28_adj_2205), 
         .D(recv_buffer[87]), .Z(n39_adj_2202)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(recv_buffer[90]), .B(n38_adj_2206), .C(n32_adj_2207), 
         .D(recv_buffer[85]), .Z(n40_adj_2203)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(recv_buffer[75]), .B(recv_buffer[82]), .C(recv_buffer[92]), 
         .D(recv_buffer[86]), .Z(n36_adj_2204)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(recv_buffer[76]), .B(recv_buffer[77]), .Z(n28_adj_2205)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(recv_buffer[83]), .B(n34_adj_2208), .C(n24_adj_2209), 
         .D(recv_buffer[91]), .Z(n38_adj_2206)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(recv_buffer[81]), .B(recv_buffer[78]), .C(recv_buffer[89]), 
         .Z(n32_adj_2207)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(recv_buffer[95]), .B(recv_buffer[94]), .C(recv_buffer[84]), 
         .D(recv_buffer[79]), .Z(n34_adj_2208)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(recv_buffer[93]), .B(recv_buffer[80]), .Z(n24_adj_2209)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i2_4_lut_adj_140 (.A(n3388), .B(n3364), .C(n39_adj_2210), .D(n40_adj_2211), 
         .Z(enable_m2_N_635)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_140.init = 16'h8880;
    LUT4 i18_4_lut_adj_141 (.A(recv_buffer[67]), .B(n36_adj_2212), .C(n28_adj_2213), 
         .D(recv_buffer[66]), .Z(n39_adj_2210)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_141.init = 16'hfffe;
    LUT4 i19_4_lut_adj_142 (.A(recv_buffer[69]), .B(n38_adj_2214), .C(n32_adj_2215), 
         .D(recv_buffer[64]), .Z(n40_adj_2211)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_142.init = 16'hfffe;
    LUT4 i15_4_lut_adj_143 (.A(recv_buffer[54]), .B(recv_buffer[61]), .C(recv_buffer[71]), 
         .D(recv_buffer[65]), .Z(n36_adj_2212)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_143.init = 16'hfffe;
    LUT4 i7_2_lut_adj_144 (.A(recv_buffer[55]), .B(recv_buffer[56]), .Z(n28_adj_2213)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_144.init = 16'heeee;
    LUT4 i17_4_lut_adj_145 (.A(recv_buffer[62]), .B(n34_adj_2216), .C(n24_adj_2217), 
         .D(recv_buffer[70]), .Z(n38_adj_2214)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_145.init = 16'hfffe;
    LUT4 i11_3_lut_adj_146 (.A(recv_buffer[60]), .B(recv_buffer[57]), .C(recv_buffer[68]), 
         .Z(n32_adj_2215)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_146.init = 16'hfefe;
    LUT4 i13_4_lut_adj_147 (.A(recv_buffer[74]), .B(recv_buffer[73]), .C(recv_buffer[63]), 
         .D(recv_buffer[58]), .Z(n34_adj_2216)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_147.init = 16'hfffe;
    LUT4 i3_2_lut_adj_148 (.A(recv_buffer[72]), .B(recv_buffer[59]), .Z(n24_adj_2217)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_148.init = 16'heeee;
    LUT4 i2_4_lut_adj_149 (.A(n3436), .B(n3412), .C(n39_adj_2218), .D(n40_adj_2219), 
         .Z(enable_m3_N_642)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_149.init = 16'h8880;
    LUT4 i18_4_lut_adj_150 (.A(recv_buffer[46]), .B(n36_adj_2220), .C(n28_adj_2221), 
         .D(recv_buffer[45]), .Z(n39_adj_2218)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_150.init = 16'hfffe;
    LUT4 i19_4_lut_adj_151 (.A(recv_buffer[48]), .B(n38_adj_2222), .C(n32_adj_2223), 
         .D(recv_buffer[43]), .Z(n40_adj_2219)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_151.init = 16'hfffe;
    FD1P3AX send_buffer_i0_i1 (.D(send_buffer_95__N_346[1]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i1.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i2 (.D(send_buffer_95__N_346[2]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i3 (.D(send_buffer_95__N_346[3]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i4 (.D(send_buffer_95__N_346[4]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i4.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i5 (.D(send_buffer_95__N_346[5]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i5.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i6 (.D(send_buffer_95__N_346[6]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i7 (.D(send_buffer_95__N_346[7]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i8 (.D(send_buffer_95__N_346[8]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i8.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i9 (.D(send_buffer_95__N_346[9]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i9.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i10 (.D(send_buffer_95__N_346[10]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i10.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i11 (.D(send_buffer_95__N_346[11]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i11.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i12 (.D(send_buffer_95__N_346[12]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i12.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i13 (.D(send_buffer_95__N_346[13]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i13.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i14 (.D(send_buffer_95__N_346[14]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i14.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i15 (.D(send_buffer_95__N_346[15]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i15.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i16 (.D(send_buffer_95__N_346[16]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i16.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i17 (.D(send_buffer_95__N_346[17]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i17.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i18 (.D(send_buffer_95__N_346[18]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i18.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i19 (.D(send_buffer_95__N_346[19]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i19.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i20 (.D(send_buffer_95__N_346[20]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i20.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i21 (.D(send_buffer_95__N_346[21]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i21.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i22 (.D(send_buffer_95__N_346[22]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i22.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i23 (.D(send_buffer_95__N_346[23]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i23.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i24 (.D(send_buffer_95__N_346[24]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i24.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i25 (.D(send_buffer_95__N_346[25]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i25.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i26 (.D(send_buffer_95__N_346[26]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i26.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i27 (.D(send_buffer_95__N_346[27]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i27.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i28 (.D(send_buffer_95__N_346[28]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i28.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i29 (.D(send_buffer_95__N_346[29]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i29.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i30 (.D(send_buffer_95__N_346[30]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i30.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i31 (.D(send_buffer_95__N_346[31]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i31.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i32 (.D(send_buffer_95__N_346[32]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i32.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i33 (.D(send_buffer_95__N_346[33]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i33.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i34 (.D(send_buffer_95__N_346[34]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i34.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i35 (.D(send_buffer_95__N_346[35]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i35.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i36 (.D(send_buffer_95__N_346[36]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i36.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i37 (.D(send_buffer_95__N_346[37]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i37.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i38 (.D(send_buffer_95__N_346[38]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i38.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i39 (.D(send_buffer_95__N_346[39]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i39.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i40 (.D(send_buffer_95__N_346[40]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i40.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i41 (.D(send_buffer_95__N_346[41]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i41.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i42 (.D(send_buffer_95__N_346[42]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i42.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i43 (.D(send_buffer_95__N_346[43]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i43.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i44 (.D(send_buffer_95__N_346[44]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i44.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i45 (.D(send_buffer_95__N_346[45]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i45.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i46 (.D(send_buffer_95__N_346[46]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i46.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i47 (.D(send_buffer_95__N_346[47]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i47.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i48 (.D(send_buffer_95__N_346[48]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i48.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i49 (.D(send_buffer_95__N_346[49]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i49.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i50 (.D(send_buffer_95__N_346[50]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i50.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i51 (.D(send_buffer_95__N_346[51]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i51.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i52 (.D(send_buffer_95__N_346[52]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i52.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i53 (.D(send_buffer_95__N_346[53]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i53.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i54 (.D(send_buffer_95__N_346[54]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i54.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i55 (.D(send_buffer_95__N_346[55]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i55.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i56 (.D(send_buffer_95__N_346[56]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i56.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i57 (.D(send_buffer_95__N_346[57]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i57.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i58 (.D(send_buffer_95__N_346[58]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i58.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i59 (.D(send_buffer_95__N_346[59]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i59.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i60 (.D(send_buffer_95__N_346[60]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i60.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i61 (.D(send_buffer_95__N_346[61]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i61.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i62 (.D(send_buffer_95__N_346[62]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i62.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i63 (.D(send_buffer_95__N_346[63]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i63.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i64 (.D(send_buffer_95__N_346[64]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i64.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i65 (.D(send_buffer_95__N_346[65]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i65.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i66 (.D(send_buffer_95__N_346[66]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i66.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i67 (.D(send_buffer_95__N_346[67]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i67.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i68 (.D(send_buffer_95__N_346[68]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i68.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i69 (.D(send_buffer_95__N_346[69]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i69.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i70 (.D(send_buffer_95__N_346[70]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i70.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i71 (.D(send_buffer_95__N_346[71]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i71.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i72 (.D(send_buffer_95__N_346[72]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i72.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i73 (.D(send_buffer_95__N_346[73]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i73.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i74 (.D(send_buffer_95__N_346[74]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i74.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i75 (.D(send_buffer_95__N_346[75]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i75.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i76 (.D(send_buffer_95__N_346[76]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i76.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i77 (.D(send_buffer_95__N_346[77]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i77.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i78 (.D(send_buffer_95__N_346[78]), .SP(clkout_c_enable_172), 
            .CK(clkout_c), .Q(send_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i78.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i79 (.D(send_buffer_95__N_346[79]), .SP(clkout_c_enable_173), 
            .CK(clkout_c), .Q(send_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i79.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i80 (.D(send_buffer_95__N_346[80]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i80.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i81 (.D(send_buffer_95__N_346[81]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i81.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i82 (.D(send_buffer_95__N_346[82]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i82.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i83 (.D(send_buffer_95__N_346[83]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i83.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i84 (.D(send_buffer_95__N_346[84]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i84.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i85 (.D(send_buffer_95__N_346[85]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i85.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i86 (.D(send_buffer_95__N_346[86]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i86.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i87 (.D(send_buffer_95__N_346[87]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i87.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i88 (.D(send_buffer_95__N_346[88]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i88.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i89 (.D(send_buffer_95__N_346[89]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i89.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i90 (.D(send_buffer_95__N_346[90]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i90.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i91 (.D(send_buffer_95__N_346[91]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i91.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i92 (.D(send_buffer_95__N_346[92]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i92.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i93 (.D(send_buffer_95__N_346[93]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i93.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i94 (.D(\send_buffer_95__N_346[94] ), .SP(rst), 
            .CK(clkout_c), .Q(\send_buffer[94] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i94.GSR = "DISABLED";
    LUT4 i15_4_lut_adj_152 (.A(recv_buffer[33]), .B(recv_buffer[40]), .C(recv_buffer[50]), 
         .D(recv_buffer[44]), .Z(n36_adj_2220)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_152.init = 16'hfffe;
    LUT4 i7_2_lut_adj_153 (.A(recv_buffer[34]), .B(recv_buffer[35]), .Z(n28_adj_2221)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_153.init = 16'heeee;
    LUT4 i2_4_lut_adj_154 (.A(n3484), .B(n3460), .C(n39_adj_2224), .D(n40_adj_2225), 
         .Z(enable_m4_N_649)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_154.init = 16'h8880;
    LUT4 i17_4_lut_adj_155 (.A(recv_buffer[41]), .B(n34_adj_2226), .C(n24_adj_2227), 
         .D(recv_buffer[49]), .Z(n38_adj_2222)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_155.init = 16'hfffe;
    LUT4 i18_4_lut_adj_156 (.A(recv_buffer[25]), .B(n36_adj_2228), .C(n28_adj_2229), 
         .D(recv_buffer[24]), .Z(n39_adj_2224)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_156.init = 16'hfffe;
    LUT4 i19_4_lut_adj_157 (.A(recv_buffer[27]), .B(n38_adj_2230), .C(n32_adj_2231), 
         .D(recv_buffer[22]), .Z(n40_adj_2225)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_157.init = 16'hfffe;
    LUT4 i11_3_lut_adj_158 (.A(recv_buffer[39]), .B(recv_buffer[36]), .C(recv_buffer[47]), 
         .Z(n32_adj_2223)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_158.init = 16'hfefe;
    LUT4 i13_4_lut_adj_159 (.A(recv_buffer[53]), .B(recv_buffer[52]), .C(recv_buffer[42]), 
         .D(recv_buffer[37]), .Z(n34_adj_2226)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_159.init = 16'hfffe;
    LUT4 i3_2_lut_adj_160 (.A(recv_buffer[51]), .B(recv_buffer[38]), .Z(n24_adj_2227)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_160.init = 16'heeee;
    CCU2D add_15010_2 (.A0(recv_buffer[59]), .B0(recv_buffer[58]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[60]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18272));
    defparam add_15010_2.INIT0 = 16'h7000;
    defparam add_15010_2.INIT1 = 16'h5aaa;
    defparam add_15010_2.INJECT1_0 = "NO";
    defparam add_15010_2.INJECT1_1 = "NO";
    CCU2D add_15011_21 (.A0(recv_buffer[74]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18271), .S1(n3364));
    defparam add_15011_21.INIT0 = 16'h5555;
    defparam add_15011_21.INIT1 = 16'h0000;
    defparam add_15011_21.INJECT1_0 = "NO";
    defparam add_15011_21.INJECT1_1 = "NO";
    LUT4 mux_51_i2_3_lut_4_lut_else_4_lut (.A(CSlatched), .B(send_buffer[1]), 
         .C(CSold), .Z(n22086)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i2_3_lut_4_lut_else_4_lut.init = 16'hdcdc;
    LUT4 i15_4_lut_adj_161 (.A(n169[0]), .B(recv_buffer[19]), .C(recv_buffer[29]), 
         .D(recv_buffer[23]), .Z(n36_adj_2228)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_161.init = 16'hfffe;
    LUT4 CSlatched_I_0_1_lut (.A(CSlatched), .Z(CSlatched_N_664)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam CSlatched_I_0_1_lut.init = 16'h5555;
    LUT4 i3_4_lut (.A(SCKold), .B(n22100), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_94)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut.init = 16'h0400;
    CCU2D add_15011_19 (.A0(recv_buffer[72]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[73]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18270), .COUT(n18271));
    defparam add_15011_19.INIT0 = 16'hf555;
    defparam add_15011_19.INIT1 = 16'hf555;
    defparam add_15011_19.INJECT1_0 = "NO";
    defparam add_15011_19.INJECT1_1 = "NO";
    LUT4 i7_2_lut_adj_162 (.A(recv_buffer[13]), .B(recv_buffer[14]), .Z(n28_adj_2229)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_162.init = 16'heeee;
    LUT4 i2_3_lut_rep_371 (.A(CSlatched), .B(CSold), .C(n22100), .Z(clkout_c_enable_254)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i2_3_lut_rep_371.init = 16'h8080;
    LUT4 i11648_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22100), .D(enable_m1_N_627), 
         .Z(n14202)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11648_2_lut_4_lut.init = 16'h0080;
    LUT4 i11628_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22100), .D(enable_m2_N_635), 
         .Z(n14182)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11628_2_lut_4_lut.init = 16'h0080;
    LUT4 i11608_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22100), .D(enable_m3_N_642), 
         .Z(n14162)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11608_2_lut_4_lut.init = 16'h0080;
    LUT4 i11588_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22100), .D(enable_m4_N_649), 
         .Z(n14142)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11588_2_lut_4_lut.init = 16'h0080;
    CCU2D add_15011_17 (.A0(recv_buffer[70]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[71]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18269), .COUT(n18270));
    defparam add_15011_17.INIT0 = 16'hf555;
    defparam add_15011_17.INIT1 = 16'hf555;
    defparam add_15011_17.INJECT1_0 = "NO";
    defparam add_15011_17.INJECT1_1 = "NO";
    CCU2D add_15011_15 (.A0(recv_buffer[68]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[69]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18268), .COUT(n18269));
    defparam add_15011_15.INIT0 = 16'hf555;
    defparam add_15011_15.INIT1 = 16'hf555;
    defparam add_15011_15.INJECT1_0 = "NO";
    defparam add_15011_15.INJECT1_1 = "NO";
    CCU2D add_15011_13 (.A0(recv_buffer[66]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[67]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18267), .COUT(n18268));
    defparam add_15011_13.INIT0 = 16'hf555;
    defparam add_15011_13.INIT1 = 16'h0aaa;
    defparam add_15011_13.INJECT1_0 = "NO";
    defparam add_15011_13.INJECT1_1 = "NO";
    LUT4 i17_4_lut_adj_163 (.A(recv_buffer[20]), .B(n34_adj_2232), .C(n24_adj_2233), 
         .D(recv_buffer[28]), .Z(n38_adj_2230)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_163.init = 16'hfffe;
    LUT4 CSold_I_0_2_lut_rep_373 (.A(CSold), .B(CSlatched), .Z(n21354)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam CSold_I_0_2_lut_rep_373.init = 16'h2222;
    LUT4 mux_9_i76_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[0] ), 
         .D(send_buffer[75]), .Z(MISOb_N_666[75])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i76_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i84_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[8] ), 
         .D(send_buffer[83]), .Z(MISOb_N_666[83])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i84_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i85_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[9] ), 
         .D(send_buffer[84]), .Z(MISOb_N_666[84])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i85_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13072_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[19] ), 
         .D(send_buffer[73]), .Z(MISOb_N_666[73])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13072_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i86_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[10] ), 
         .D(send_buffer[85]), .Z(MISOb_N_666[85])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i86_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11_3_lut_adj_164 (.A(recv_buffer[18]), .B(recv_buffer[15]), .C(recv_buffer[26]), 
         .Z(n32_adj_2231)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_164.init = 16'hfefe;
    LUT4 i13_4_lut_adj_165 (.A(recv_buffer[32]), .B(recv_buffer[31]), .C(recv_buffer[21]), 
         .D(recv_buffer[16]), .Z(n34_adj_2232)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_165.init = 16'hfffe;
    LUT4 i3_2_lut_adj_166 (.A(recv_buffer[30]), .B(recv_buffer[17]), .Z(n24_adj_2233)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_166.init = 16'heeee;
    LUT4 i13132_2_lut_3_lut (.A(n22098), .B(CSlatched), .C(send_buffer[74]), 
         .Z(MISOb_N_666[74])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13132_2_lut_3_lut.init = 16'hd0d0;
    CCU2D add_15011_11 (.A0(recv_buffer[64]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[65]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18266), .COUT(n18267));
    defparam add_15011_11.INIT0 = 16'h0aaa;
    defparam add_15011_11.INIT1 = 16'hf555;
    defparam add_15011_11.INJECT1_0 = "NO";
    defparam add_15011_11.INJECT1_1 = "NO";
    CCU2D add_15011_9 (.A0(recv_buffer[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18265), .COUT(n18266));
    defparam add_15011_9.INIT0 = 16'h0aaa;
    defparam add_15011_9.INIT1 = 16'h0aaa;
    defparam add_15011_9.INJECT1_0 = "NO";
    defparam add_15011_9.INJECT1_1 = "NO";
    LUT4 mux_9_i82_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[6] ), 
         .D(send_buffer[81]), .Z(MISOb_N_666[81])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i82_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i83_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[7] ), 
         .D(send_buffer[82]), .Z(MISOb_N_666[82])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i83_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i80_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[4] ), 
         .D(send_buffer[79]), .Z(MISOb_N_666[79])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i80_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i78_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[2] ), 
         .D(send_buffer[77]), .Z(MISOb_N_666[77])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i78_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i77_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[1] ), 
         .D(send_buffer[76]), .Z(MISOb_N_666[76])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i77_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i79_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[3] ), 
         .D(send_buffer[78]), .Z(MISOb_N_666[78])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i79_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i81_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[5] ), 
         .D(send_buffer[80]), .Z(MISOb_N_666[80])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i81_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i87_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[11] ), 
         .D(send_buffer[86]), .Z(MISOb_N_666[86])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i87_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i88_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[12] ), 
         .D(send_buffer[87]), .Z(MISOb_N_666[87])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i88_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i89_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[13] ), 
         .D(send_buffer[88]), .Z(MISOb_N_666[88])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i89_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i90_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[14] ), 
         .D(send_buffer[89]), .Z(MISOb_N_666[89])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i90_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i91_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[15] ), 
         .D(send_buffer[90]), .Z(MISOb_N_666[90])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i91_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i92_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[16] ), 
         .D(send_buffer[91]), .Z(MISOb_N_666[91])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i92_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i93_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[17] ), 
         .D(send_buffer[92]), .Z(MISOb_N_666[92])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i93_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i94_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[18] ), 
         .D(send_buffer[93]), .Z(MISOb_N_666[93])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i94_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i21_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[8] ), 
         .D(send_buffer[20]), .Z(MISOb_N_666[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[7] ), 
         .D(send_buffer[19]), .Z(MISOb_N_666[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i20_3_lut_4_lut.init = 16'hfd20;
    PFUMX i17311 (.BLUT(n21289), .ALUT(n21288), .C0(n22100), .Z(MISO_N_670));
    LUT4 mux_9_i23_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[10] ), 
         .D(send_buffer[22]), .Z(MISOb_N_666[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i22_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[9] ), 
         .D(send_buffer[21]), .Z(MISOb_N_666[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i24_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[11] ), 
         .D(send_buffer[23]), .Z(MISOb_N_666[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i24_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15011_7 (.A0(recv_buffer[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18264), .COUT(n18265));
    defparam add_15011_7.INIT0 = 16'hf555;
    defparam add_15011_7.INIT1 = 16'hf555;
    defparam add_15011_7.INJECT1_0 = "NO";
    defparam add_15011_7.INJECT1_1 = "NO";
    CCU2D add_15011_5 (.A0(recv_buffer[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18263), .COUT(n18264));
    defparam add_15011_5.INIT0 = 16'h0aaa;
    defparam add_15011_5.INIT1 = 16'hf555;
    defparam add_15011_5.INJECT1_0 = "NO";
    defparam add_15011_5.INJECT1_1 = "NO";
    LUT4 mux_9_i25_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[12] ), 
         .D(send_buffer[24]), .Z(MISOb_N_666[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i25_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15011_3 (.A0(recv_buffer[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18262), .COUT(n18263));
    defparam add_15011_3.INIT0 = 16'hf555;
    defparam add_15011_3.INIT1 = 16'hf555;
    defparam add_15011_3.INJECT1_0 = "NO";
    defparam add_15011_3.INJECT1_1 = "NO";
    LUT4 mux_9_i26_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[13] ), 
         .D(send_buffer[25]), .Z(MISOb_N_666[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i26_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15011_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[54]), .B1(recv_buffer[55]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18262));
    defparam add_15011_1.INIT0 = 16'hF000;
    defparam add_15011_1.INIT1 = 16'ha666;
    defparam add_15011_1.INJECT1_0 = "NO";
    defparam add_15011_1.INJECT1_1 = "NO";
    LUT4 mux_9_i27_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[14] ), 
         .D(send_buffer[26]), .Z(MISOb_N_666[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i27_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15012_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18261), 
          .S0(n3436));
    defparam add_15012_cout.INIT0 = 16'h0000;
    defparam add_15012_cout.INIT1 = 16'h0000;
    defparam add_15012_cout.INJECT1_0 = "NO";
    defparam add_15012_cout.INJECT1_1 = "NO";
    LUT4 mux_9_i28_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[15] ), 
         .D(send_buffer[27]), .Z(MISOb_N_666[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i29_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[16] ), 
         .D(send_buffer[28]), .Z(MISOb_N_666[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i30_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[17] ), 
         .D(send_buffer[29]), .Z(MISOb_N_666[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i31_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[18] ), 
         .D(send_buffer[30]), .Z(MISOb_N_666[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i31_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13074_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[19] ), 
         .D(send_buffer[31]), .Z(MISOb_N_666[31])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13074_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(enable_m4), 
         .D(send_buffer[8]), .Z(MISOb_N_666[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13234_2_lut_3_lut (.A(n22098), .B(CSlatched), .C(send_buffer[7]), 
         .Z(MISOb_N_666[7])) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13234_2_lut_3_lut.init = 16'hf2f2;
    CCU2D add_15012_16 (.A0(recv_buffer[52]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[53]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18260), .COUT(n18261));
    defparam add_15012_16.INIT0 = 16'h5aaa;
    defparam add_15012_16.INIT1 = 16'h0aaa;
    defparam add_15012_16.INJECT1_0 = "NO";
    defparam add_15012_16.INJECT1_1 = "NO";
    CCU2D add_15012_14 (.A0(recv_buffer[50]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[51]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18259), .COUT(n18260));
    defparam add_15012_14.INIT0 = 16'h5aaa;
    defparam add_15012_14.INIT1 = 16'h5aaa;
    defparam add_15012_14.INJECT1_0 = "NO";
    defparam add_15012_14.INJECT1_1 = "NO";
    CCU2D add_14993_21 (.A0(recv_buffer[95]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18102), .S1(n3316));
    defparam add_14993_21.INIT0 = 16'h5555;
    defparam add_14993_21.INIT1 = 16'h0000;
    defparam add_14993_21.INJECT1_0 = "NO";
    defparam add_14993_21.INJECT1_1 = "NO";
    CCU2D add_15012_12 (.A0(recv_buffer[48]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[49]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18258), .COUT(n18259));
    defparam add_15012_12.INIT0 = 16'h5aaa;
    defparam add_15012_12.INIT1 = 16'h5aaa;
    defparam add_15012_12.INJECT1_0 = "NO";
    defparam add_15012_12.INJECT1_1 = "NO";
    CCU2D add_14993_19 (.A0(recv_buffer[93]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[94]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18101), .COUT(n18102));
    defparam add_14993_19.INIT0 = 16'hf555;
    defparam add_14993_19.INIT1 = 16'hf555;
    defparam add_14993_19.INJECT1_0 = "NO";
    defparam add_14993_19.INJECT1_1 = "NO";
    CCU2D add_14993_17 (.A0(recv_buffer[91]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[92]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18100), .COUT(n18101));
    defparam add_14993_17.INIT0 = 16'hf555;
    defparam add_14993_17.INIT1 = 16'hf555;
    defparam add_14993_17.INJECT1_0 = "NO";
    defparam add_14993_17.INJECT1_1 = "NO";
    CCU2D add_15012_10 (.A0(recv_buffer[46]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[47]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18257), .COUT(n18258));
    defparam add_15012_10.INIT0 = 16'h5555;
    defparam add_15012_10.INIT1 = 16'h5aaa;
    defparam add_15012_10.INJECT1_0 = "NO";
    defparam add_15012_10.INJECT1_1 = "NO";
    CCU2D add_14993_15 (.A0(recv_buffer[89]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[90]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18099), .COUT(n18100));
    defparam add_14993_15.INIT0 = 16'hf555;
    defparam add_14993_15.INIT1 = 16'hf555;
    defparam add_14993_15.INJECT1_0 = "NO";
    defparam add_14993_15.INJECT1_1 = "NO";
    CCU2D add_15012_8 (.A0(recv_buffer[44]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[45]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18256), .COUT(n18257));
    defparam add_15012_8.INIT0 = 16'h5aaa;
    defparam add_15012_8.INIT1 = 16'h5aaa;
    defparam add_15012_8.INJECT1_0 = "NO";
    defparam add_15012_8.INJECT1_1 = "NO";
    CCU2D add_15012_6 (.A0(recv_buffer[42]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[43]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18255), .COUT(n18256));
    defparam add_15012_6.INIT0 = 16'h5555;
    defparam add_15012_6.INIT1 = 16'h5555;
    defparam add_15012_6.INJECT1_0 = "NO";
    defparam add_15012_6.INJECT1_1 = "NO";
    CCU2D add_15012_4 (.A0(recv_buffer[40]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[41]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18254), .COUT(n18255));
    defparam add_15012_4.INIT0 = 16'h5aaa;
    defparam add_15012_4.INIT1 = 16'h5555;
    defparam add_15012_4.INJECT1_0 = "NO";
    defparam add_15012_4.INJECT1_1 = "NO";
    CCU2D add_14993_13 (.A0(recv_buffer[87]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[88]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18098), .COUT(n18099));
    defparam add_14993_13.INIT0 = 16'hf555;
    defparam add_14993_13.INIT1 = 16'h0aaa;
    defparam add_14993_13.INJECT1_0 = "NO";
    defparam add_14993_13.INJECT1_1 = "NO";
    CCU2D add_15012_2 (.A0(recv_buffer[38]), .B0(recv_buffer[37]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[39]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18254));
    defparam add_15012_2.INIT0 = 16'h7000;
    defparam add_15012_2.INIT1 = 16'h5aaa;
    defparam add_15012_2.INJECT1_0 = "NO";
    defparam add_15012_2.INJECT1_1 = "NO";
    LUT4 i13196_2_lut_3_lut (.A(n22098), .B(CSlatched), .C(send_buffer[32]), 
         .Z(MISOb_N_666[32])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13196_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_9_i34_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[0] ), 
         .D(send_buffer[33]), .Z(MISOb_N_666[33])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i34_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i35_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[1] ), 
         .D(send_buffer[34]), .Z(MISOb_N_666[34])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i35_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i36_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[2] ), 
         .D(send_buffer[35]), .Z(MISOb_N_666[35])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i36_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i37_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[3] ), 
         .D(send_buffer[36]), .Z(MISOb_N_666[36])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i37_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i38_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[4] ), 
         .D(send_buffer[37]), .Z(MISOb_N_666[37])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i38_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i39_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[5] ), 
         .D(send_buffer[38]), .Z(MISOb_N_666[38])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i39_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i40_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[6] ), 
         .D(send_buffer[39]), .Z(MISOb_N_666[39])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i40_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i41_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[7] ), 
         .D(send_buffer[40]), .Z(MISOb_N_666[40])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i41_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_14993_11 (.A0(recv_buffer[85]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[86]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18097), .COUT(n18098));
    defparam add_14993_11.INIT0 = 16'h0aaa;
    defparam add_14993_11.INIT1 = 16'hf555;
    defparam add_14993_11.INJECT1_0 = "NO";
    defparam add_14993_11.INJECT1_1 = "NO";
    LUT4 mux_9_i42_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[8] ), 
         .D(send_buffer[41]), .Z(MISOb_N_666[41])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i42_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_14993_9 (.A0(recv_buffer[83]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[84]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18096), .COUT(n18097));
    defparam add_14993_9.INIT0 = 16'h0aaa;
    defparam add_14993_9.INIT1 = 16'h0aaa;
    defparam add_14993_9.INJECT1_0 = "NO";
    defparam add_14993_9.INJECT1_1 = "NO";
    CCU2D add_14993_7 (.A0(recv_buffer[81]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[82]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18095), .COUT(n18096));
    defparam add_14993_7.INIT0 = 16'hf555;
    defparam add_14993_7.INIT1 = 16'hf555;
    defparam add_14993_7.INJECT1_0 = "NO";
    defparam add_14993_7.INJECT1_1 = "NO";
    CCU2D add_14993_5 (.A0(recv_buffer[79]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[80]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18094), .COUT(n18095));
    defparam add_14993_5.INIT0 = 16'h0aaa;
    defparam add_14993_5.INIT1 = 16'hf555;
    defparam add_14993_5.INJECT1_0 = "NO";
    defparam add_14993_5.INJECT1_1 = "NO";
    CCU2D add_14993_3 (.A0(recv_buffer[77]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[78]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18093), .COUT(n18094));
    defparam add_14993_3.INIT0 = 16'hf555;
    defparam add_14993_3.INIT1 = 16'hf555;
    defparam add_14993_3.INJECT1_0 = "NO";
    defparam add_14993_3.INJECT1_1 = "NO";
    CCU2D add_14993_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[75]), .B1(recv_buffer[76]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18093));
    defparam add_14993_1.INIT0 = 16'hF000;
    defparam add_14993_1.INIT1 = 16'ha666;
    defparam add_14993_1.INJECT1_0 = "NO";
    defparam add_14993_1.INJECT1_1 = "NO";
    LUT4 mux_9_i43_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[9] ), 
         .D(send_buffer[42]), .Z(MISOb_N_666[42])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i43_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i44_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[10] ), 
         .D(send_buffer[43]), .Z(MISOb_N_666[43])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i44_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i45_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[11] ), 
         .D(send_buffer[44]), .Z(MISOb_N_666[44])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i45_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX speed_set_m2_i0_i0 (.D(recv_buffer[54]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i0.GSR = "DISABLED";
    LUT4 mux_9_i46_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[12] ), 
         .D(send_buffer[45]), .Z(MISOb_N_666[45])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i46_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i47_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[13] ), 
         .D(send_buffer[46]), .Z(MISOb_N_666[46])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i47_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i48_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[14] ), 
         .D(send_buffer[47]), .Z(MISOb_N_666[47])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i48_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX speed_set_m1_i0_i0 (.D(recv_buffer[75]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i0.GSR = "DISABLED";
    LUT4 mux_9_i49_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[15] ), 
         .D(send_buffer[48]), .Z(MISOb_N_666[48])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i49_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i50_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[16] ), 
         .D(send_buffer[49]), .Z(MISOb_N_666[49])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i50_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i51_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[17] ), 
         .D(send_buffer[50]), .Z(MISOb_N_666[50])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i51_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i52_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[18] ), 
         .D(send_buffer[51]), .Z(MISOb_N_666[51])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i52_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(enable_m2), 
         .D(send_buffer[10]), .Z(MISOb_N_666[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(enable_m3), 
         .D(send_buffer[9]), .Z(MISOb_N_666[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13073_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m3[19] ), 
         .D(send_buffer[52]), .Z(MISOb_N_666[52])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13073_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13178_2_lut_3_lut (.A(n22098), .B(CSlatched), .C(send_buffer[53]), 
         .Z(MISOb_N_666[53])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13178_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_9_i55_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[0] ), 
         .D(send_buffer[54]), .Z(MISOb_N_666[54])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i55_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i56_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[1] ), 
         .D(send_buffer[55]), .Z(MISOb_N_666[55])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i56_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i57_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[2] ), 
         .D(send_buffer[56]), .Z(MISOb_N_666[56])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i57_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i58_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[3] ), 
         .D(send_buffer[57]), .Z(MISOb_N_666[57])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i58_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i59_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[4] ), 
         .D(send_buffer[58]), .Z(MISOb_N_666[58])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i59_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i60_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[5] ), 
         .D(send_buffer[59]), .Z(MISOb_N_666[59])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i60_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i61_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[6] ), 
         .D(send_buffer[60]), .Z(MISOb_N_666[60])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i61_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i62_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[7] ), 
         .D(send_buffer[61]), .Z(MISOb_N_666[61])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i62_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i63_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[8] ), 
         .D(send_buffer[62]), .Z(MISOb_N_666[62])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i63_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i64_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[9] ), 
         .D(send_buffer[63]), .Z(MISOb_N_666[63])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i64_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i65_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[10] ), 
         .D(send_buffer[64]), .Z(MISOb_N_666[64])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i65_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i66_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[11] ), 
         .D(send_buffer[65]), .Z(MISOb_N_666[65])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i66_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i67_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[12] ), 
         .D(send_buffer[66]), .Z(MISOb_N_666[66])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i67_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i68_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[13] ), 
         .D(send_buffer[67]), .Z(MISOb_N_666[67])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i68_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i69_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[14] ), 
         .D(send_buffer[68]), .Z(MISOb_N_666[68])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i69_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i70_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[15] ), 
         .D(send_buffer[69]), .Z(MISOb_N_666[69])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i70_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i71_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[16] ), 
         .D(send_buffer[70]), .Z(MISOb_N_666[70])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i71_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i72_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[17] ), 
         .D(send_buffer[71]), .Z(MISOb_N_666[71])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i72_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i73_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m2[18] ), 
         .D(send_buffer[72]), .Z(MISOb_N_666[72])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i73_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(enable_m1), 
         .D(send_buffer[11]), .Z(MISOb_N_666[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[0] ), 
         .D(send_buffer[12]), .Z(MISOb_N_666[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13238_2_lut_3_lut (.A(n22098), .B(CSlatched), .C(send_buffer[3]), 
         .Z(MISOb_N_666[3])) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13238_2_lut_3_lut.init = 16'hf2f2;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[1] ), 
         .D(send_buffer[13]), .Z(MISOb_N_666[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13061_3_lut_rep_354_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m1[19] ), 
         .D(\send_buffer[94] ), .Z(n21335)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13061_3_lut_rep_354_4_lut.init = 16'hfd20;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[2] ), 
         .D(send_buffer[14]), .Z(MISOb_N_666[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13237_2_lut_3_lut (.A(n22098), .B(CSlatched), .C(send_buffer[4]), 
         .Z(MISOb_N_666[4])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13237_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[3] ), 
         .D(send_buffer[15]), .Z(MISOb_N_666[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13236_2_lut_3_lut (.A(CSold), .B(CSlatched), .C(send_buffer[5]), 
         .Z(MISOb_N_666[5])) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13236_2_lut_3_lut.init = 16'hf2f2;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[4] ), 
         .D(send_buffer[16]), .Z(MISOb_N_666[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[5] ), 
         .D(send_buffer[17]), .Z(MISOb_N_666[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13235_2_lut_3_lut (.A(CSold), .B(CSlatched), .C(send_buffer[6]), 
         .Z(MISOb_N_666[6])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam i13235_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n22098), .B(CSlatched), .C(\speed_avg_m4[6] ), 
         .D(send_buffer[18]), .Z(MISOb_N_666[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[7:42])
    defparam mux_9_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 SCKold_I_0_2_lut_rep_374 (.A(SCKold), .B(SCKlatched), .Z(n21355)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(193[8:45])
    defparam SCKold_I_0_2_lut_rep_374.init = 16'h2222;
    LUT4 i131_2_lut_rep_355_3_lut (.A(SCKold), .B(SCKlatched), .C(CSlatched), 
         .Z(n21336)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(193[8:45])
    defparam i131_2_lut_rep_355_3_lut.init = 16'h0202;
    LUT4 i2716_1_lut (.A(MISO_N_625), .Z(n5132)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    defparam i2716_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_379 (.A(enable_m4), .B(free_m4), .Z(n21360)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_379.init = 16'h2222;
    LUT4 i17179_3_lut_4_lut (.A(enable_m4), .B(free_m4), .C(hallsense_m4[2]), 
         .D(hallsense_m4[0]), .Z(n19415)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17179_3_lut_4_lut.init = 16'hfddf;
    FD1P3IX speed_set_m4_i0_i12 (.D(recv_buffer[24]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_384 (.A(enable_m3), .B(free_m3), .Z(n21365)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_384.init = 16'h2222;
    LUT4 i17169_3_lut_4_lut (.A(enable_m3), .B(free_m3), .C(hallsense_m3[2]), 
         .D(hallsense_m3[0]), .Z(n19427)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17169_3_lut_4_lut.init = 16'hfddf;
    LUT4 i1_2_lut_rep_389 (.A(enable_m2), .B(free_m2), .Z(n21370)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_389.init = 16'h2222;
    LUT4 i17159_3_lut_4_lut (.A(enable_m2), .B(free_m2), .C(hallsense_m2[2]), 
         .D(hallsense_m2[0]), .Z(n19411)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17159_3_lut_4_lut.init = 16'hfddf;
    LUT4 i1_2_lut_rep_393 (.A(enable_m1), .B(free_m1), .Z(n21374)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i1_2_lut_rep_393.init = 16'h2222;
    LUT4 i17149_3_lut_4_lut (.A(enable_m1), .B(free_m1), .C(hallsense_m1[2]), 
         .D(hallsense_m1[0]), .Z(n19421)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i17149_3_lut_4_lut.init = 16'hfddf;
    FD1P3JX speed_set_m4_i0_i13 (.D(recv_buffer[25]), .SP(clkout_c_enable_254), 
            .PD(n14142), .CK(clkout_c), .Q(speed_set_m4[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i14 (.D(recv_buffer[26]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i1 (.D(recv_buffer[76]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i2 (.D(recv_buffer[77]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i3 (.D(recv_buffer[78]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i4 (.D(recv_buffer[79]), .SP(clkout_c_enable_254), 
            .PD(n14202), .CK(clkout_c), .Q(speed_set_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i5 (.D(recv_buffer[80]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i6 (.D(recv_buffer[81]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i7 (.D(recv_buffer[82]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i8 (.D(recv_buffer[83]), .SP(clkout_c_enable_254), 
            .PD(n14202), .CK(clkout_c), .Q(speed_set_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i9 (.D(recv_buffer[84]), .SP(clkout_c_enable_254), 
            .PD(n14202), .CK(clkout_c), .Q(speed_set_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i10 (.D(recv_buffer[85]), .SP(clkout_c_enable_254), 
            .PD(n14202), .CK(clkout_c), .Q(speed_set_m1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i11 (.D(recv_buffer[86]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i12 (.D(recv_buffer[87]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i13 (.D(recv_buffer[88]), .SP(clkout_c_enable_254), 
            .PD(n14202), .CK(clkout_c), .Q(speed_set_m1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i14 (.D(recv_buffer[89]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i15 (.D(recv_buffer[90]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i16 (.D(recv_buffer[91]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i17 (.D(recv_buffer[92]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i18 (.D(recv_buffer[93]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i19 (.D(recv_buffer[94]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i20 (.D(recv_buffer[95]), .SP(clkout_c_enable_254), 
            .CD(n14202), .CK(clkout_c), .Q(speed_set_m1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i1 (.D(recv_buffer[55]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i2 (.D(recv_buffer[56]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i3 (.D(recv_buffer[57]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i4 (.D(recv_buffer[58]), .SP(clkout_c_enable_254), 
            .PD(n14182), .CK(clkout_c), .Q(speed_set_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i5 (.D(recv_buffer[59]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i6 (.D(recv_buffer[60]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i7 (.D(recv_buffer[61]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i8 (.D(recv_buffer[62]), .SP(clkout_c_enable_254), 
            .PD(n14182), .CK(clkout_c), .Q(speed_set_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i9 (.D(recv_buffer[63]), .SP(clkout_c_enable_254), 
            .PD(n14182), .CK(clkout_c), .Q(speed_set_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i10 (.D(recv_buffer[64]), .SP(clkout_c_enable_254), 
            .PD(n14182), .CK(clkout_c), .Q(speed_set_m2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i11 (.D(recv_buffer[65]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i12 (.D(recv_buffer[66]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i13 (.D(recv_buffer[67]), .SP(clkout_c_enable_254), 
            .PD(n14182), .CK(clkout_c), .Q(speed_set_m2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i14 (.D(recv_buffer[68]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i15 (.D(recv_buffer[69]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i16 (.D(recv_buffer[70]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i17 (.D(recv_buffer[71]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i18 (.D(recv_buffer[72]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i19 (.D(recv_buffer[73]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i20 (.D(recv_buffer[74]), .SP(clkout_c_enable_254), 
            .CD(n14182), .CK(clkout_c), .Q(speed_set_m2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i1 (.D(recv_buffer[34]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i2 (.D(recv_buffer[35]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i3 (.D(recv_buffer[36]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i4 (.D(recv_buffer[37]), .SP(clkout_c_enable_254), 
            .PD(n14162), .CK(clkout_c), .Q(speed_set_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i5 (.D(recv_buffer[38]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i6 (.D(recv_buffer[39]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i7 (.D(recv_buffer[40]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i8 (.D(recv_buffer[41]), .SP(clkout_c_enable_254), 
            .PD(n14162), .CK(clkout_c), .Q(speed_set_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i9 (.D(recv_buffer[42]), .SP(clkout_c_enable_254), 
            .PD(n14162), .CK(clkout_c), .Q(speed_set_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i10 (.D(recv_buffer[43]), .SP(clkout_c_enable_254), 
            .PD(n14162), .CK(clkout_c), .Q(speed_set_m3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i11 (.D(recv_buffer[44]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i12 (.D(recv_buffer[45]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i12.GSR = "DISABLED";
    CCU2D add_15007_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18307), 
          .S0(n3484));
    defparam add_15007_cout.INIT0 = 16'h0000;
    defparam add_15007_cout.INIT1 = 16'h0000;
    defparam add_15007_cout.INJECT1_0 = "NO";
    defparam add_15007_cout.INJECT1_1 = "NO";
    FD1P3JX speed_set_m3_i0_i13 (.D(recv_buffer[46]), .SP(clkout_c_enable_254), 
            .PD(n14162), .CK(clkout_c), .Q(speed_set_m3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i14 (.D(recv_buffer[47]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i15 (.D(recv_buffer[48]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i16 (.D(recv_buffer[49]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i17 (.D(recv_buffer[50]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i18 (.D(recv_buffer[51]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i19 (.D(recv_buffer[52]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i20 (.D(recv_buffer[53]), .SP(clkout_c_enable_254), 
            .CD(n14162), .CK(clkout_c), .Q(speed_set_m3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i1 (.D(recv_buffer[13]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i2 (.D(recv_buffer[14]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i3 (.D(recv_buffer[15]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i4 (.D(recv_buffer[16]), .SP(clkout_c_enable_254), 
            .PD(n14142), .CK(clkout_c), .Q(speed_set_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i5 (.D(recv_buffer[17]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i6 (.D(recv_buffer[18]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i7 (.D(recv_buffer[19]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i8 (.D(recv_buffer[20]), .SP(clkout_c_enable_254), 
            .PD(n14142), .CK(clkout_c), .Q(speed_set_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i9 (.D(recv_buffer[21]), .SP(clkout_c_enable_254), 
            .PD(n14142), .CK(clkout_c), .Q(speed_set_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i10 (.D(recv_buffer[22]), .SP(clkout_c_enable_254), 
            .PD(n14142), .CK(clkout_c), .Q(speed_set_m4[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i10.GSR = "DISABLED";
    CCU2D add_15007_16 (.A0(recv_buffer[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[32]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18306), .COUT(n18307));
    defparam add_15007_16.INIT0 = 16'h5aaa;
    defparam add_15007_16.INIT1 = 16'h0aaa;
    defparam add_15007_16.INJECT1_0 = "NO";
    defparam add_15007_16.INJECT1_1 = "NO";
    CCU2D add_14992_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18072), 
          .S0(n3340));
    defparam add_14992_cout.INIT0 = 16'h0000;
    defparam add_14992_cout.INIT1 = 16'h0000;
    defparam add_14992_cout.INJECT1_0 = "NO";
    defparam add_14992_cout.INJECT1_1 = "NO";
    CCU2D add_15007_14 (.A0(recv_buffer[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18305), .COUT(n18306));
    defparam add_15007_14.INIT0 = 16'h5aaa;
    defparam add_15007_14.INIT1 = 16'h5aaa;
    defparam add_15007_14.INJECT1_0 = "NO";
    defparam add_15007_14.INJECT1_1 = "NO";
    CCU2D add_15007_12 (.A0(recv_buffer[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18304), .COUT(n18305));
    defparam add_15007_12.INIT0 = 16'h5aaa;
    defparam add_15007_12.INIT1 = 16'h5aaa;
    defparam add_15007_12.INJECT1_0 = "NO";
    defparam add_15007_12.INJECT1_1 = "NO";
    CCU2D add_14992_16 (.A0(recv_buffer[94]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[95]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18071), .COUT(n18072));
    defparam add_14992_16.INIT0 = 16'h5aaa;
    defparam add_14992_16.INIT1 = 16'h0aaa;
    defparam add_14992_16.INJECT1_0 = "NO";
    defparam add_14992_16.INJECT1_1 = "NO";
    LUT4 mux_51_i3_3_lut_4_lut_then_4_lut (.A(CSlatched), .B(send_buffer[2]), 
         .C(CSold), .D(send_buffer[3]), .Z(n22091)) /* synthesis lut_function=(A (B)+!A (C+(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i3_3_lut_4_lut_then_4_lut.init = 16'hddd8;
    CCU2D add_14992_14 (.A0(recv_buffer[92]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[93]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18070), .COUT(n18071));
    defparam add_14992_14.INIT0 = 16'h5aaa;
    defparam add_14992_14.INIT1 = 16'h5aaa;
    defparam add_14992_14.INJECT1_0 = "NO";
    defparam add_14992_14.INJECT1_1 = "NO";
    CCU2D add_14992_12 (.A0(recv_buffer[90]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[91]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18069), .COUT(n18070));
    defparam add_14992_12.INIT0 = 16'h5aaa;
    defparam add_14992_12.INIT1 = 16'h5aaa;
    defparam add_14992_12.INJECT1_0 = "NO";
    defparam add_14992_12.INJECT1_1 = "NO";
    CCU2D add_14992_10 (.A0(recv_buffer[88]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[89]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18068), .COUT(n18069));
    defparam add_14992_10.INIT0 = 16'h5555;
    defparam add_14992_10.INIT1 = 16'h5aaa;
    defparam add_14992_10.INJECT1_0 = "NO";
    defparam add_14992_10.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i15 (.D(recv_buffer[27]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i15.GSR = "DISABLED";
    CCU2D add_15007_10 (.A0(recv_buffer[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18303), .COUT(n18304));
    defparam add_15007_10.INIT0 = 16'h5555;
    defparam add_15007_10.INIT1 = 16'h5aaa;
    defparam add_15007_10.INJECT1_0 = "NO";
    defparam add_15007_10.INJECT1_1 = "NO";
    CCU2D add_15007_8 (.A0(recv_buffer[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18302), .COUT(n18303));
    defparam add_15007_8.INIT0 = 16'h5aaa;
    defparam add_15007_8.INIT1 = 16'h5aaa;
    defparam add_15007_8.INJECT1_0 = "NO";
    defparam add_15007_8.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i16 (.D(recv_buffer[28]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i16.GSR = "DISABLED";
    CCU2D add_15007_6 (.A0(recv_buffer[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18301), .COUT(n18302));
    defparam add_15007_6.INIT0 = 16'h5555;
    defparam add_15007_6.INIT1 = 16'h5555;
    defparam add_15007_6.INJECT1_0 = "NO";
    defparam add_15007_6.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i17 (.D(recv_buffer[29]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i17.GSR = "DISABLED";
    LUT4 mux_51_i3_3_lut_4_lut_else_4_lut (.A(CSlatched), .B(send_buffer[2]), 
         .C(CSold), .Z(n22090)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(192[3] 206[10])
    defparam mux_51_i3_3_lut_4_lut_else_4_lut.init = 16'h8c8c;
    CCU2D add_15007_4 (.A0(recv_buffer[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18300), .COUT(n18301));
    defparam add_15007_4.INIT0 = 16'h5aaa;
    defparam add_15007_4.INIT1 = 16'h5555;
    defparam add_15007_4.INJECT1_0 = "NO";
    defparam add_15007_4.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i11 (.D(recv_buffer[23]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i18 (.D(recv_buffer[30]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i19 (.D(recv_buffer[31]), .SP(clkout_c_enable_254), 
            .CD(n14142), .CK(clkout_c), .Q(speed_set_m4[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=307, LSE_RLINE=307 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i19.GSR = "DISABLED";
    CCU2D add_14992_8 (.A0(recv_buffer[86]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[87]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18067), .COUT(n18068));
    defparam add_14992_8.INIT0 = 16'h5aaa;
    defparam add_14992_8.INIT1 = 16'h5aaa;
    defparam add_14992_8.INJECT1_0 = "NO";
    defparam add_14992_8.INJECT1_1 = "NO";
    CCU2D add_15007_2 (.A0(recv_buffer[17]), .B0(recv_buffer[16]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18300));
    defparam add_15007_2.INIT0 = 16'h7000;
    defparam add_15007_2.INIT1 = 16'h5aaa;
    defparam add_15007_2.INJECT1_0 = "NO";
    defparam add_15007_2.INJECT1_1 = "NO";
    CCU2D add_15008_21 (.A0(recv_buffer[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18299), .S1(n3460));
    defparam add_15008_21.INIT0 = 16'h5555;
    defparam add_15008_21.INIT1 = 16'h0000;
    defparam add_15008_21.INJECT1_0 = "NO";
    defparam add_15008_21.INJECT1_1 = "NO";
    CCU2D add_14992_6 (.A0(recv_buffer[84]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[85]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18066), .COUT(n18067));
    defparam add_14992_6.INIT0 = 16'h5555;
    defparam add_14992_6.INIT1 = 16'h5555;
    defparam add_14992_6.INJECT1_0 = "NO";
    defparam add_14992_6.INJECT1_1 = "NO";
    CCU2D add_15008_19 (.A0(recv_buffer[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18298), .COUT(n18299));
    defparam add_15008_19.INIT0 = 16'hf555;
    defparam add_15008_19.INIT1 = 16'hf555;
    defparam add_15008_19.INJECT1_0 = "NO";
    defparam add_15008_19.INJECT1_1 = "NO";
    CCU2D add_15008_17 (.A0(recv_buffer[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18297), .COUT(n18298));
    defparam add_15008_17.INIT0 = 16'hf555;
    defparam add_15008_17.INIT1 = 16'hf555;
    defparam add_15008_17.INJECT1_0 = "NO";
    defparam add_15008_17.INJECT1_1 = "NO";
    CCU2D add_15008_15 (.A0(recv_buffer[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18296), .COUT(n18297));
    defparam add_15008_15.INIT0 = 16'hf555;
    defparam add_15008_15.INIT1 = 16'hf555;
    defparam add_15008_15.INJECT1_0 = "NO";
    defparam add_15008_15.INJECT1_1 = "NO";
    CCU2D add_14992_4 (.A0(recv_buffer[82]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[83]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18065), .COUT(n18066));
    defparam add_14992_4.INIT0 = 16'h5aaa;
    defparam add_14992_4.INIT1 = 16'h5555;
    defparam add_14992_4.INJECT1_0 = "NO";
    defparam add_14992_4.INJECT1_1 = "NO";
    CCU2D add_15008_13 (.A0(recv_buffer[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18295), .COUT(n18296));
    defparam add_15008_13.INIT0 = 16'hf555;
    defparam add_15008_13.INIT1 = 16'h0aaa;
    defparam add_15008_13.INJECT1_0 = "NO";
    defparam add_15008_13.INJECT1_1 = "NO";
    CCU2D add_15008_11 (.A0(recv_buffer[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18294), .COUT(n18295));
    defparam add_15008_11.INIT0 = 16'h0aaa;
    defparam add_15008_11.INIT1 = 16'hf555;
    defparam add_15008_11.INJECT1_0 = "NO";
    defparam add_15008_11.INJECT1_1 = "NO";
    CCU2D add_15008_9 (.A0(recv_buffer[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18293), .COUT(n18294));
    defparam add_15008_9.INIT0 = 16'h0aaa;
    defparam add_15008_9.INIT1 = 16'h0aaa;
    defparam add_15008_9.INJECT1_0 = "NO";
    defparam add_15008_9.INJECT1_1 = "NO";
    CCU2D add_15008_7 (.A0(recv_buffer[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18292), .COUT(n18293));
    defparam add_15008_7.INIT0 = 16'hf555;
    defparam add_15008_7.INIT1 = 16'hf555;
    defparam add_15008_7.INJECT1_0 = "NO";
    defparam add_15008_7.INJECT1_1 = "NO";
    CCU2D add_15008_5 (.A0(recv_buffer[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18291), .COUT(n18292));
    defparam add_15008_5.INIT0 = 16'h0aaa;
    defparam add_15008_5.INIT1 = 16'hf555;
    defparam add_15008_5.INJECT1_0 = "NO";
    defparam add_15008_5.INJECT1_1 = "NO";
    CCU2D add_15008_3 (.A0(recv_buffer[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18290), .COUT(n18291));
    defparam add_15008_3.INIT0 = 16'hf555;
    defparam add_15008_3.INIT1 = 16'hf555;
    defparam add_15008_3.INJECT1_0 = "NO";
    defparam add_15008_3.INJECT1_1 = "NO";
    CCU2D add_14992_2 (.A0(recv_buffer[80]), .B0(recv_buffer[79]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[81]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18065));
    defparam add_14992_2.INIT0 = 16'h7000;
    defparam add_14992_2.INIT1 = 16'h5aaa;
    defparam add_14992_2.INJECT1_0 = "NO";
    defparam add_14992_2.INJECT1_1 = "NO";
    CCU2D add_15008_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n169[0]), .B1(recv_buffer[13]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18290));
    defparam add_15008_1.INIT0 = 16'hF000;
    defparam add_15008_1.INIT1 = 16'ha666;
    defparam add_15008_1.INJECT1_0 = "NO";
    defparam add_15008_1.INJECT1_1 = "NO";
    CCU2D add_15009_21 (.A0(recv_buffer[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18289), .S1(n3412));
    defparam add_15009_21.INIT0 = 16'h5555;
    defparam add_15009_21.INIT1 = 16'h0000;
    defparam add_15009_21.INJECT1_0 = "NO";
    defparam add_15009_21.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U0
//

module PWMGENERATOR_U0 (PWM_m3, pwm_clk, free_m3, rst, PWMdut_m3, 
            GND_net, hallsense_m3, n21363, enable_m3, n3124, n21366, 
            n3088);
    output PWM_m3;
    input pwm_clk;
    output free_m3;
    input rst;
    input [9:0]PWMdut_m3;
    input GND_net;
    input [2:0]hallsense_m3;
    output n21363;
    input enable_m3;
    output n3124;
    output n21366;
    output n3088;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_1982, free_N_1994, n10, n7, n10_adj_2200, n11407, 
        n9, n3871, n18207;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    wire [9:0]n45;
    
    wire n19794, n6, n14138, n19740, n18206, n18205, n18204, n18203, 
        n14, n10_adj_2201, n18159, n18158, n18157, n18156, n18155;
    
    FD1S3AX PWM_20 (.D(PWM_N_1982), .CK(pwm_clk), .Q(PWM_m3)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1994), .SP(rst), .CK(pwm_clk), .Q(free_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(PWMdut_m3[5]), .B(PWMdut_m3[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_2200), .B(PWMdut_m3[9]), .C(PWMdut_m3[8]), 
         .D(PWMdut_m3[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2292_3_lut (.A(n11407), .B(PWMdut_m3[4]), .C(PWMdut_m3[3]), 
         .Z(n10_adj_2200)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2292_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1796_1_lut (.A(n3871), .Z(PWM_N_1982)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1796_1_lut.init = 16'h5555;
    CCU2D cnt_2084_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18207), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2084_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2084_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2084_add_4_11.INJECT1_1 = "NO";
    LUT4 i17118_4_lut (.A(cnt[2]), .B(n19794), .C(cnt[1]), .D(n6), .Z(n14138)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17118_4_lut.init = 16'h0004;
    LUT4 i16403_3_lut (.A(cnt[6]), .B(n19740), .C(cnt[8]), .Z(n19794)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16403_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[4]), .B(cnt[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i16351_4_lut (.A(cnt[7]), .B(cnt[5]), .C(cnt[9]), .D(cnt[3]), 
         .Z(n19740)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16351_4_lut.init = 16'h8000;
    CCU2D cnt_2084_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18206), 
          .COUT(n18207), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2084_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2084_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2084_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2084_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18205), 
          .COUT(n18206), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2084_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2084_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2084_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2084_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18204), 
          .COUT(n18205), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2084_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2084_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2084_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2084_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18203), 
          .COUT(n18204), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2084_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2084_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2084_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2084_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18203), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2084_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2084_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2084_add_4_1.INJECT1_1 = "NO";
    LUT4 i17090_4_lut (.A(PWMdut_m3[5]), .B(n14), .C(n10_adj_2201), .D(PWMdut_m3[8]), 
         .Z(free_N_1994)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17090_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m3[9]), .B(PWMdut_m3[3]), .C(PWMdut_m3[4]), 
         .D(n11407), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m3[6]), .B(PWMdut_m3[7]), .Z(n10_adj_2201)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_132 (.A(PWMdut_m3[2]), .B(PWMdut_m3[1]), .C(PWMdut_m3[0]), 
         .Z(n11407)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_132.init = 16'hfefe;
    LUT4 i1620_3_lut_rep_382 (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .Z(n21363)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1620_3_lut_rep_382.init = 16'h1414;
    LUT4 i17165_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[0]), .C(hallsense_m3[1]), 
         .D(enable_m3), .Z(n3124)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17165_2_lut_4_lut.init = 16'hebff;
    LUT4 i1590_3_lut_rep_385 (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .Z(n21366)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1590_3_lut_rep_385.init = 16'h1414;
    LUT4 i17162_2_lut_4_lut (.A(free_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .D(enable_m3), .Z(n3088)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17162_2_lut_4_lut.init = 16'hebff;
    CCU2D sub_1794_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m3[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18159), .S1(n3871));
    defparam sub_1794_add_2_11.INIT0 = 16'h5999;
    defparam sub_1794_add_2_11.INIT1 = 16'h0000;
    defparam sub_1794_add_2_11.INJECT1_0 = "NO";
    defparam sub_1794_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_9 (.A0(PWMdut_m3[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m3[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18158), 
          .COUT(n18159));
    defparam sub_1794_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1794_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1794_add_2_9.INJECT1_0 = "NO";
    defparam sub_1794_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_7 (.A0(PWMdut_m3[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m3[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18157), 
          .COUT(n18158));
    defparam sub_1794_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1794_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1794_add_2_7.INJECT1_0 = "NO";
    defparam sub_1794_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_5 (.A0(PWMdut_m3[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m3[4]), .C1(n9), .D1(n10), .CIN(n18156), 
          .COUT(n18157));
    defparam sub_1794_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1794_add_2_5.INIT1 = 16'h5999;
    defparam sub_1794_add_2_5.INJECT1_0 = "NO";
    defparam sub_1794_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m3[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m3[2]), .C1(n9), .D1(n10), .CIN(n18155), 
          .COUT(n18156));
    defparam sub_1794_add_2_3.INIT0 = 16'h5999;
    defparam sub_1794_add_2_3.INIT1 = 16'h5999;
    defparam sub_1794_add_2_3.INJECT1_0 = "NO";
    defparam sub_1794_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1794_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m3[0]), .C1(n9), .D1(n10), 
          .COUT(n18155));
    defparam sub_1794_add_2_1.INIT0 = 16'h0000;
    defparam sub_1794_add_2_1.INIT1 = 16'h5999;
    defparam sub_1794_add_2_1.INJECT1_0 = "NO";
    defparam sub_1794_add_2_1.INJECT1_1 = "NO";
    FD1S3IX cnt_2084__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14138), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i0.GSR = "ENABLED";
    FD1S3IX cnt_2084__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14138), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i1.GSR = "ENABLED";
    FD1S3IX cnt_2084__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14138), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i2.GSR = "ENABLED";
    FD1S3IX cnt_2084__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14138), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i3.GSR = "ENABLED";
    FD1S3IX cnt_2084__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14138), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i4.GSR = "ENABLED";
    FD1S3IX cnt_2084__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14138), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i5.GSR = "ENABLED";
    FD1S3IX cnt_2084__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14138), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i6.GSR = "ENABLED";
    FD1S3IX cnt_2084__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14138), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i7.GSR = "ENABLED";
    FD1S3IX cnt_2084__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14138), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i8.GSR = "ENABLED";
    FD1S3IX cnt_2084__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14138), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2084__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U1
//

module PWMGENERATOR_U1 (PWMdut_m2, GND_net, PWM_m2, pwm_clk, free_m2, 
            rst, hallsense_m2, n21369, enable_m2, n3016, n21371, 
            n2980);
    input [9:0]PWMdut_m2;
    input GND_net;
    output PWM_m2;
    input pwm_clk;
    output free_m2;
    input rst;
    input [2:0]hallsense_m2;
    output n21369;
    input enable_m2;
    output n3016;
    output n21371;
    output n2980;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire n9, n18212;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    wire [9:0]n45;
    
    wire PWM_N_1982, n18211, n18210, n18209, free_N_1994, n3858, 
        n18208, n19796, n6, n14139, n19744, n14, n10, n11405, 
        n18164, n18163, n7, n18162, n18161, n10_adj_2198, n18160, 
        n10_adj_2199;
    
    LUT4 i3_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D cnt_2083_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18212), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2083_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2083_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2083_add_4_11.INJECT1_1 = "NO";
    FD1S3AX PWM_20 (.D(PWM_N_1982), .CK(pwm_clk), .Q(PWM_m2)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    CCU2D cnt_2083_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18211), 
          .COUT(n18212), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2083_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2083_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2083_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2083_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18210), 
          .COUT(n18211), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2083_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2083_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2083_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2083_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18209), 
          .COUT(n18210), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2083_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2083_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2083_add_4_5.INJECT1_1 = "NO";
    FD1P3AX free_19 (.D(free_N_1994), .SP(rst), .CK(pwm_clk), .Q(free_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i1794_1_lut (.A(n3858), .Z(PWM_N_1982)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1794_1_lut.init = 16'h5555;
    CCU2D cnt_2083_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18208), 
          .COUT(n18209), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2083_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2083_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2083_add_4_3.INJECT1_1 = "NO";
    LUT4 i17121_4_lut (.A(cnt[0]), .B(n19796), .C(cnt[2]), .D(n6), .Z(n14139)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17121_4_lut.init = 16'h0004;
    LUT4 i16405_3_lut (.A(cnt[7]), .B(n19744), .C(cnt[3]), .Z(n19796)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16405_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i16355_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n19744)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16355_4_lut.init = 16'h8000;
    CCU2D cnt_2083_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18208), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2083_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2083_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2083_add_4_1.INJECT1_1 = "NO";
    LUT4 i17096_4_lut (.A(PWMdut_m2[5]), .B(n14), .C(n10), .D(PWMdut_m2[8]), 
         .Z(free_N_1994)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17096_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m2[9]), .B(PWMdut_m2[3]), .C(PWMdut_m2[4]), 
         .D(n11405), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m2[6]), .B(PWMdut_m2[7]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(PWMdut_m2[2]), .B(PWMdut_m2[1]), .C(PWMdut_m2[0]), 
         .Z(n11405)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut.init = 16'hfefe;
    CCU2D sub_1792_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m2[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18164), .S1(n3858));
    defparam sub_1792_add_2_11.INIT0 = 16'h5999;
    defparam sub_1792_add_2_11.INIT1 = 16'h0000;
    defparam sub_1792_add_2_11.INJECT1_0 = "NO";
    defparam sub_1792_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_9 (.A0(PWMdut_m2[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m2[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18163), 
          .COUT(n18164));
    defparam sub_1792_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1792_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1792_add_2_9.INJECT1_0 = "NO";
    defparam sub_1792_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_7 (.A0(PWMdut_m2[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m2[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18162), 
          .COUT(n18163));
    defparam sub_1792_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1792_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1792_add_2_7.INJECT1_0 = "NO";
    defparam sub_1792_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_5 (.A0(PWMdut_m2[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m2[4]), .C1(n9), .D1(n10_adj_2198), 
          .CIN(n18161), .COUT(n18162));
    defparam sub_1792_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1792_add_2_5.INIT1 = 16'h5999;
    defparam sub_1792_add_2_5.INJECT1_0 = "NO";
    defparam sub_1792_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m2[1]), .C0(n9), .D0(n10_adj_2198), 
          .A1(cnt[2]), .B1(PWMdut_m2[2]), .C1(n9), .D1(n10_adj_2198), 
          .CIN(n18160), .COUT(n18161));
    defparam sub_1792_add_2_3.INIT0 = 16'h5999;
    defparam sub_1792_add_2_3.INIT1 = 16'h5999;
    defparam sub_1792_add_2_3.INJECT1_0 = "NO";
    defparam sub_1792_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1792_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m2[0]), .C1(n9), .D1(n10_adj_2198), 
          .COUT(n18160));
    defparam sub_1792_add_2_1.INIT0 = 16'h0000;
    defparam sub_1792_add_2_1.INIT1 = 16'h5999;
    defparam sub_1792_add_2_1.INJECT1_0 = "NO";
    defparam sub_1792_add_2_1.INJECT1_1 = "NO";
    LUT4 i1530_3_lut_rep_388 (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .Z(n21369)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1530_3_lut_rep_388.init = 16'h1414;
    LUT4 i17155_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[0]), .C(hallsense_m2[1]), 
         .D(enable_m2), .Z(n3016)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17155_2_lut_4_lut.init = 16'hebff;
    LUT4 i1500_3_lut_rep_390 (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .Z(n21371)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1500_3_lut_rep_390.init = 16'h1414;
    LUT4 i17152_2_lut_4_lut (.A(free_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .D(enable_m2), .Z(n2980)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17152_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2083__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14139), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i0.GSR = "ENABLED";
    LUT4 i2_3_lut_adj_131 (.A(PWMdut_m2[5]), .B(PWMdut_m2[6]), .C(n10_adj_2198), 
         .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_adj_131.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_2199), .B(PWMdut_m2[9]), .C(PWMdut_m2[8]), 
         .D(PWMdut_m2[7]), .Z(n10_adj_2198)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2282_3_lut (.A(n11405), .B(PWMdut_m2[4]), .C(PWMdut_m2[3]), 
         .Z(n10_adj_2199)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2282_3_lut.init = 16'hecec;
    FD1S3IX cnt_2083__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14139), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i1.GSR = "ENABLED";
    FD1S3IX cnt_2083__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14139), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i2.GSR = "ENABLED";
    FD1S3IX cnt_2083__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14139), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i3.GSR = "ENABLED";
    FD1S3IX cnt_2083__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14139), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i4.GSR = "ENABLED";
    FD1S3IX cnt_2083__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14139), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i5.GSR = "ENABLED";
    FD1S3IX cnt_2083__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14139), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i6.GSR = "ENABLED";
    FD1S3IX cnt_2083__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14139), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i7.GSR = "ENABLED";
    FD1S3IX cnt_2083__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14139), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i8.GSR = "ENABLED";
    FD1S3IX cnt_2083__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14139), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2083__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U2
//

module PWMGENERATOR_U2 (GND_net, PWM_m1, pwm_clk, free_m1, rst, PWMdut_m1, 
            hallsense_m1, n21373, enable_m1, n2908, n21375, n2872);
    input GND_net;
    output PWM_m1;
    input pwm_clk;
    output free_m1;
    input rst;
    input [9:0]PWMdut_m1;
    input [2:0]hallsense_m1;
    output n21373;
    input enable_m1;
    output n2908;
    output n21375;
    output n2872;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire n18217;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    wire [9:0]n45;
    
    wire n18216, n18215, n18214, n18213, PWM_N_1982, n3845, free_N_1994, 
        n17, n16, n14140, n10, n7, n10_adj_2196, n11403, n9, 
        n14, n10_adj_2197, n18169, n18168, n18167, n18166, n18165;
    
    CCU2D cnt_2082_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18217), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2082_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2082_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2082_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2082_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18216), 
          .COUT(n18217), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2082_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2082_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2082_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2082_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18215), 
          .COUT(n18216), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2082_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2082_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2082_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2082_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18214), 
          .COUT(n18215), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2082_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2082_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2082_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2082_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18213), 
          .COUT(n18214), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2082_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2082_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2082_add_4_3.INJECT1_1 = "NO";
    FD1S3AX PWM_20 (.D(PWM_N_1982), .CK(pwm_clk), .Q(PWM_m1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    CCU2D cnt_2082_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18213), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2082_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2082_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2082_add_4_1.INJECT1_1 = "NO";
    LUT4 i1792_1_lut (.A(n3845), .Z(PWM_N_1982)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1792_1_lut.init = 16'h5555;
    FD1P3AX free_19 (.D(free_N_1994), .SP(rst), .CK(pwm_clk), .Q(free_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i17124_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n14140)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17124_4_lut.init = 16'h0400;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i6_4_lut (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut.init = 16'hffef;
    LUT4 i2_3_lut (.A(PWMdut_m1[5]), .B(PWMdut_m1[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_2196), .B(PWMdut_m1[9]), .C(PWMdut_m1[8]), 
         .D(PWMdut_m1[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2272_3_lut (.A(n11403), .B(PWMdut_m1[4]), .C(PWMdut_m1[3]), 
         .Z(n10_adj_2196)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2272_3_lut.init = 16'hecec;
    LUT4 i3_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i17099_4_lut (.A(PWMdut_m1[5]), .B(n14), .C(n10_adj_2197), .D(PWMdut_m1[8]), 
         .Z(free_N_1994)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17099_4_lut.init = 16'h0001;
    LUT4 i6_4_lut_adj_129 (.A(PWMdut_m1[9]), .B(PWMdut_m1[3]), .C(PWMdut_m1[4]), 
         .D(n11403), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut_adj_129.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[7]), .Z(n10_adj_2197)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_130 (.A(PWMdut_m1[2]), .B(PWMdut_m1[1]), .C(PWMdut_m1[0]), 
         .Z(n11403)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_130.init = 16'hfefe;
    CCU2D sub_1790_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m1[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18169), .S1(n3845));
    defparam sub_1790_add_2_11.INIT0 = 16'h5999;
    defparam sub_1790_add_2_11.INIT1 = 16'h0000;
    defparam sub_1790_add_2_11.INJECT1_0 = "NO";
    defparam sub_1790_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_9 (.A0(PWMdut_m1[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m1[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18168), 
          .COUT(n18169));
    defparam sub_1790_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1790_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1790_add_2_9.INJECT1_0 = "NO";
    defparam sub_1790_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_7 (.A0(PWMdut_m1[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m1[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18167), 
          .COUT(n18168));
    defparam sub_1790_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1790_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1790_add_2_7.INJECT1_0 = "NO";
    defparam sub_1790_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_5 (.A0(PWMdut_m1[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m1[4]), .C1(n9), .D1(n10), .CIN(n18166), 
          .COUT(n18167));
    defparam sub_1790_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1790_add_2_5.INIT1 = 16'h5999;
    defparam sub_1790_add_2_5.INJECT1_0 = "NO";
    defparam sub_1790_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m1[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m1[2]), .C1(n9), .D1(n10), .CIN(n18165), 
          .COUT(n18166));
    defparam sub_1790_add_2_3.INIT0 = 16'h5999;
    defparam sub_1790_add_2_3.INIT1 = 16'h5999;
    defparam sub_1790_add_2_3.INJECT1_0 = "NO";
    defparam sub_1790_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1790_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m1[0]), .C1(n9), .D1(n10), 
          .COUT(n18165));
    defparam sub_1790_add_2_1.INIT0 = 16'h0000;
    defparam sub_1790_add_2_1.INIT1 = 16'h5999;
    defparam sub_1790_add_2_1.INJECT1_0 = "NO";
    defparam sub_1790_add_2_1.INJECT1_1 = "NO";
    LUT4 i1440_3_lut_rep_392 (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .Z(n21373)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1440_3_lut_rep_392.init = 16'h1414;
    LUT4 i17145_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[0]), .C(hallsense_m1[1]), 
         .D(enable_m1), .Z(n2908)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17145_2_lut_4_lut.init = 16'hebff;
    LUT4 i1410_3_lut_rep_394 (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .Z(n21375)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1410_3_lut_rep_394.init = 16'h1414;
    LUT4 i17142_2_lut_4_lut (.A(free_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .D(enable_m1), .Z(n2872)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17142_2_lut_4_lut.init = 16'hebff;
    FD1S3IX cnt_2082__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14140), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i0.GSR = "ENABLED";
    FD1S3IX cnt_2082__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14140), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i1.GSR = "ENABLED";
    FD1S3IX cnt_2082__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14140), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i2.GSR = "ENABLED";
    FD1S3IX cnt_2082__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14140), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i3.GSR = "ENABLED";
    FD1S3IX cnt_2082__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14140), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i4.GSR = "ENABLED";
    FD1S3IX cnt_2082__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14140), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i5.GSR = "ENABLED";
    FD1S3IX cnt_2082__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14140), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i6.GSR = "ENABLED";
    FD1S3IX cnt_2082__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14140), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i7.GSR = "ENABLED";
    FD1S3IX cnt_2082__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14140), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i8.GSR = "ENABLED";
    FD1S3IX cnt_2082__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14140), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2082__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR
//

module PWMGENERATOR (PWM_m4, pwm_clk, free_m4, rst, PWMdut_m4, GND_net, 
            hallsense_m4, n21358, enable_m4, n3232, n21361, n3196);
    output PWM_m4;
    input pwm_clk;
    output free_m4;
    input rst;
    input [9:0]PWMdut_m4;
    input GND_net;
    input [2:0]hallsense_m4;
    output n21358;
    input enable_m4;
    output n3232;
    output n21361;
    output n3196;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_1982, free_N_1994, n3884, n10, n7, n10_adj_2194, 
        n11409, n14, n10_adj_2195, n18202;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    wire [9:0]n45;
    
    wire n18201, n18200, n18199, n18198, n9, n18154, n18153, n18152, 
        n18151, n18150, n14137, n19804, n6, n19764;
    
    FD1S3AX PWM_20 (.D(PWM_N_1982), .CK(pwm_clk), .Q(PWM_m4)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam PWM_20.GSR = "ENABLED";
    FD1P3AX free_19 (.D(free_N_1994), .SP(rst), .CK(pwm_clk), .Q(free_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam free_19.GSR = "DISABLED";
    LUT4 i1798_1_lut (.A(n3884), .Z(PWM_N_1982)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1798_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(PWMdut_m4[5]), .B(PWMdut_m4[6]), .C(n10), .Z(n7)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i3_4_lut (.A(n10_adj_2194), .B(PWMdut_m4[9]), .C(PWMdut_m4[8]), 
         .D(PWMdut_m4[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2302_3_lut (.A(n11409), .B(PWMdut_m4[4]), .C(PWMdut_m4[3]), 
         .Z(n10_adj_2194)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2302_3_lut.init = 16'hecec;
    LUT4 i17087_4_lut (.A(PWMdut_m4[5]), .B(n14), .C(n10_adj_2195), .D(PWMdut_m4[8]), 
         .Z(free_N_1994)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i17087_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(PWMdut_m4[9]), .B(PWMdut_m4[3]), .C(PWMdut_m4[4]), 
         .D(n11409), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[7]), .Z(n10_adj_2195)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_adj_128 (.A(PWMdut_m4[2]), .B(PWMdut_m4[1]), .C(PWMdut_m4[0]), 
         .Z(n11409)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut_adj_128.init = 16'hfefe;
    CCU2D cnt_2085_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18202), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2085_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2085_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2085_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2085_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18201), 
          .COUT(n18202), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2085_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2085_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2085_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2085_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18200), 
          .COUT(n18201), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2085_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2085_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2085_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2085_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18199), 
          .COUT(n18200), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2085_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2085_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2085_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2085_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18198), 
          .COUT(n18199), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2085_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2085_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2085_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2085_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18198), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2085_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2085_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2085_add_4_1.INJECT1_1 = "NO";
    LUT4 i3_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[5]), .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1710_3_lut_rep_377 (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .Z(n21358)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1710_3_lut_rep_377.init = 16'h1414;
    LUT4 i17175_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[0]), .C(hallsense_m4[1]), 
         .D(enable_m4), .Z(n3232)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17175_2_lut_4_lut.init = 16'hebff;
    LUT4 i1680_3_lut_rep_380 (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .Z(n21361)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i1680_3_lut_rep_380.init = 16'h1414;
    LUT4 i17172_2_lut_4_lut (.A(free_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .D(enable_m4), .Z(n3196)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 76[9])
    defparam i17172_2_lut_4_lut.init = 16'hebff;
    CCU2D sub_1796_add_2_11 (.A0(cnt[9]), .B0(PWMdut_m4[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18154), .S1(n3884));
    defparam sub_1796_add_2_11.INIT0 = 16'h5999;
    defparam sub_1796_add_2_11.INIT1 = 16'h0000;
    defparam sub_1796_add_2_11.INJECT1_0 = "NO";
    defparam sub_1796_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_9 (.A0(PWMdut_m4[7]), .B0(n7), .C0(cnt[7]), .D0(GND_net), 
          .A1(PWMdut_m4[8]), .B1(n7), .C1(cnt[8]), .D1(GND_net), .CIN(n18153), 
          .COUT(n18154));
    defparam sub_1796_add_2_9.INIT0 = 16'he1e1;
    defparam sub_1796_add_2_9.INIT1 = 16'he1e1;
    defparam sub_1796_add_2_9.INJECT1_0 = "NO";
    defparam sub_1796_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_7 (.A0(PWMdut_m4[5]), .B0(n7), .C0(cnt[5]), .D0(GND_net), 
          .A1(PWMdut_m4[6]), .B1(n7), .C1(cnt[6]), .D1(GND_net), .CIN(n18152), 
          .COUT(n18153));
    defparam sub_1796_add_2_7.INIT0 = 16'he1e1;
    defparam sub_1796_add_2_7.INIT1 = 16'he1e1;
    defparam sub_1796_add_2_7.INJECT1_0 = "NO";
    defparam sub_1796_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_5 (.A0(PWMdut_m4[3]), .B0(n7), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(PWMdut_m4[4]), .C1(n9), .D1(n10), .CIN(n18151), 
          .COUT(n18152));
    defparam sub_1796_add_2_5.INIT0 = 16'he1e1;
    defparam sub_1796_add_2_5.INIT1 = 16'h5999;
    defparam sub_1796_add_2_5.INJECT1_0 = "NO";
    defparam sub_1796_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_3 (.A0(cnt[1]), .B0(PWMdut_m4[1]), .C0(n9), .D0(n10), 
          .A1(cnt[2]), .B1(PWMdut_m4[2]), .C1(n9), .D1(n10), .CIN(n18150), 
          .COUT(n18151));
    defparam sub_1796_add_2_3.INIT0 = 16'h5999;
    defparam sub_1796_add_2_3.INIT1 = 16'h5999;
    defparam sub_1796_add_2_3.INJECT1_0 = "NO";
    defparam sub_1796_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1796_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(PWMdut_m4[0]), .C1(n9), .D1(n10), 
          .COUT(n18150));
    defparam sub_1796_add_2_1.INIT0 = 16'h0000;
    defparam sub_1796_add_2_1.INIT1 = 16'h5999;
    defparam sub_1796_add_2_1.INJECT1_0 = "NO";
    defparam sub_1796_add_2_1.INJECT1_1 = "NO";
    FD1S3IX cnt_2085__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14137), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i0.GSR = "ENABLED";
    LUT4 i17115_4_lut (.A(cnt[0]), .B(n19804), .C(cnt[2]), .D(n6), .Z(n14137)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(73[6:16])
    defparam i17115_4_lut.init = 16'h0004;
    LUT4 i16413_3_lut (.A(cnt[7]), .B(n19764), .C(cnt[3]), .Z(n19804)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16413_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i16375_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n19764)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16375_4_lut.init = 16'h8000;
    FD1S3IX cnt_2085__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14137), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i1.GSR = "ENABLED";
    FD1S3IX cnt_2085__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14137), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i2.GSR = "ENABLED";
    FD1S3IX cnt_2085__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14137), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i3.GSR = "ENABLED";
    FD1S3IX cnt_2085__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14137), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i4.GSR = "ENABLED";
    FD1S3IX cnt_2085__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14137), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i5.GSR = "ENABLED";
    FD1S3IX cnt_2085__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14137), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i6.GSR = "ENABLED";
    FD1S3IX cnt_2085__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14137), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i7.GSR = "ENABLED";
    FD1S3IX cnt_2085__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14137), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i8.GSR = "ENABLED";
    FD1S3IX cnt_2085__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14137), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(72[9:12])
    defparam cnt_2085__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \PID(16000000,160000000,10000000) 
//

module \PID(16000000,160000000,10000000)  (\speed_avg_m4[5] , \speed_avg_m3[5] , 
            n21328, n4322, speed_set_m2, speed_set_m3, clk_N_683, 
            n18938, speed_set_m4, \speed_avg_m4[18] , \speed_avg_m3[18] , 
            \speed_avg_m4[4] , \speed_avg_m3[4] , \speed_avg_m3[3] , \speed_avg_m2[3] , 
            \speed_avg_m4[2] , \speed_avg_m3[2] , \speed_avg_m4[1] , \speed_avg_m3[1] , 
            n7, GND_net, n4417, n4416, \speed_avg_m4[0] , \speed_avg_m3[0] , 
            \speed_avg_m4[17] , \speed_avg_m3[17] , \subOut_24__N_1177[0] , 
            speed_set_m1, \speed_avg_m4[16] , \speed_avg_m3[16] , \speed_avg_m4[15] , 
            \speed_avg_m3[15] , \speed_avg_m4[14] , \speed_avg_m3[14] , 
            \speed_avg_m4[13] , \speed_avg_m3[13] , n4419, n4418, \speed_avg_m3[12] , 
            \speed_avg_m2[12] , n22100, \speed_avg_m4[11] , \speed_avg_m3[11] , 
            \speed_avg_m4[10] , \speed_avg_m3[10] , \speed_avg_m3[9] , 
            \speed_avg_m2[9] , n4421, n4420, \speed_avg_m3[8] , \speed_avg_m2[8] , 
            n4423, n4422, \speed_avg_m3[7] , \speed_avg_m2[7] , \speed_avg_m4[6] , 
            \speed_avg_m3[6] , n4425, n4424, \speed_avg_m4[7] , \speed_avg_m1[18] , 
            \speed_avg_m2[18] , \speed_avg_m1[17] , \speed_avg_m2[17] , 
            \speed_avg_m1[16] , \speed_avg_m2[16] , \speed_avg_m1[15] , 
            \speed_avg_m2[15] , \speed_avg_m1[14] , \speed_avg_m2[14] , 
            \speed_avg_m1[13] , \speed_avg_m2[13] , \speed_avg_m1[12] , 
            \speed_avg_m1[11] , \speed_avg_m2[11] , \speed_avg_m1[10] , 
            \speed_avg_m2[10] , \speed_avg_m1[9] , \speed_avg_m1[8] , 
            \speed_avg_m1[7] , \speed_avg_m1[6] , \speed_avg_m2[6] , \speed_avg_m1[5] , 
            \speed_avg_m2[5] , \speed_avg_m1[4] , \speed_avg_m2[4] , \speed_avg_m1[3] , 
            \speed_avg_m1[2] , \speed_avg_m2[2] , \speed_avg_m1[1] , \speed_avg_m2[1] , 
            \speed_avg_m1[19] , \speed_avg_m2[19] , n5, \speed_avg_m1[0] , 
            \speed_avg_m2[0] , dir_m2, dir_m3, dir_m1, dir_m4, VCC_net, 
            \subOut_24__N_1177[1] , \subOut_24__N_1177[2] , \subOut_24__N_1177[3] , 
            \subOut_24__N_1177[4] , \subOut_24__N_1177[5] , \subOut_24__N_1177[6] , 
            \subOut_24__N_1177[7] , \subOut_24__N_1177[8] , \subOut_24__N_1177[9] , 
            \subOut_24__N_1177[10] , \subOut_24__N_1177[11] , \subOut_24__N_1177[12] , 
            \subOut_24__N_1177[13] , \subOut_24__N_1177[14] , \subOut_24__N_1177[15] , 
            \subOut_24__N_1177[16] , \subOut_24__N_1177[17] , \subOut_24__N_1177[18] , 
            \subOut_24__N_1177[19] , \subOut_24__N_1177[20] , \subOut_24__N_1177[21] , 
            \subOut_24__N_1177[24] , n4427, n4426, n4429, n4428, n4431, 
            n4430, n4433, n4432, n20284, n4435, n4434, n4436, 
            n4440, n4442, n4441, n4444, n4443, n4446, n4445, PWMdut_m4, 
            PWMdut_m3, PWMdut_m2, n4448, n4447, n4450, n4449, PWMdut_m1, 
            n4452, n4451, n4454, n4453, n4456, n4455, \speed_avg_m4[3] , 
            n4458, n4457, n4460, n4459, n4461, \speed_avg_m4[12] , 
            \speed_avg_m4[9] , \speed_avg_m4[8] , n4415, n4414);
    input \speed_avg_m4[5] ;
    input \speed_avg_m3[5] ;
    output n21328;
    output n4322;
    input [20:0]speed_set_m2;
    input [20:0]speed_set_m3;
    input clk_N_683;
    output n18938;
    input [20:0]speed_set_m4;
    input \speed_avg_m4[18] ;
    input \speed_avg_m3[18] ;
    input \speed_avg_m4[4] ;
    input \speed_avg_m3[4] ;
    input \speed_avg_m3[3] ;
    input \speed_avg_m2[3] ;
    input \speed_avg_m4[2] ;
    input \speed_avg_m3[2] ;
    input \speed_avg_m4[1] ;
    input \speed_avg_m3[1] ;
    input n7;
    input GND_net;
    output n4417;
    output n4416;
    input \speed_avg_m4[0] ;
    input \speed_avg_m3[0] ;
    input \speed_avg_m4[17] ;
    input \speed_avg_m3[17] ;
    input \subOut_24__N_1177[0] ;
    input [20:0]speed_set_m1;
    input \speed_avg_m4[16] ;
    input \speed_avg_m3[16] ;
    input \speed_avg_m4[15] ;
    input \speed_avg_m3[15] ;
    input \speed_avg_m4[14] ;
    input \speed_avg_m3[14] ;
    input \speed_avg_m4[13] ;
    input \speed_avg_m3[13] ;
    output n4419;
    output n4418;
    input \speed_avg_m3[12] ;
    input \speed_avg_m2[12] ;
    input n22100;
    input \speed_avg_m4[11] ;
    input \speed_avg_m3[11] ;
    input \speed_avg_m4[10] ;
    input \speed_avg_m3[10] ;
    input \speed_avg_m3[9] ;
    input \speed_avg_m2[9] ;
    output n4421;
    output n4420;
    input \speed_avg_m3[8] ;
    input \speed_avg_m2[8] ;
    output n4423;
    output n4422;
    input \speed_avg_m3[7] ;
    input \speed_avg_m2[7] ;
    input \speed_avg_m4[6] ;
    input \speed_avg_m3[6] ;
    output n4425;
    output n4424;
    input \speed_avg_m4[7] ;
    input \speed_avg_m1[18] ;
    input \speed_avg_m2[18] ;
    input \speed_avg_m1[17] ;
    input \speed_avg_m2[17] ;
    input \speed_avg_m1[16] ;
    input \speed_avg_m2[16] ;
    input \speed_avg_m1[15] ;
    input \speed_avg_m2[15] ;
    input \speed_avg_m1[14] ;
    input \speed_avg_m2[14] ;
    input \speed_avg_m1[13] ;
    input \speed_avg_m2[13] ;
    input \speed_avg_m1[12] ;
    input \speed_avg_m1[11] ;
    input \speed_avg_m2[11] ;
    input \speed_avg_m1[10] ;
    input \speed_avg_m2[10] ;
    input \speed_avg_m1[9] ;
    input \speed_avg_m1[8] ;
    input \speed_avg_m1[7] ;
    input \speed_avg_m1[6] ;
    input \speed_avg_m2[6] ;
    input \speed_avg_m1[5] ;
    input \speed_avg_m2[5] ;
    input \speed_avg_m1[4] ;
    input \speed_avg_m2[4] ;
    input \speed_avg_m1[3] ;
    input \speed_avg_m1[2] ;
    input \speed_avg_m2[2] ;
    input \speed_avg_m1[1] ;
    input \speed_avg_m2[1] ;
    input \speed_avg_m1[19] ;
    input \speed_avg_m2[19] ;
    output n5;
    input \speed_avg_m1[0] ;
    input \speed_avg_m2[0] ;
    output dir_m2;
    output dir_m3;
    output dir_m1;
    output dir_m4;
    input VCC_net;
    input \subOut_24__N_1177[1] ;
    input \subOut_24__N_1177[2] ;
    input \subOut_24__N_1177[3] ;
    input \subOut_24__N_1177[4] ;
    input \subOut_24__N_1177[5] ;
    input \subOut_24__N_1177[6] ;
    input \subOut_24__N_1177[7] ;
    input \subOut_24__N_1177[8] ;
    input \subOut_24__N_1177[9] ;
    input \subOut_24__N_1177[10] ;
    input \subOut_24__N_1177[11] ;
    input \subOut_24__N_1177[12] ;
    input \subOut_24__N_1177[13] ;
    input \subOut_24__N_1177[14] ;
    input \subOut_24__N_1177[15] ;
    input \subOut_24__N_1177[16] ;
    input \subOut_24__N_1177[17] ;
    input \subOut_24__N_1177[18] ;
    input \subOut_24__N_1177[19] ;
    input \subOut_24__N_1177[20] ;
    input \subOut_24__N_1177[21] ;
    input \subOut_24__N_1177[24] ;
    output n4427;
    output n4426;
    output n4429;
    output n4428;
    output n4431;
    output n4430;
    output n4433;
    output n4432;
    output n20284;
    output n4435;
    output n4434;
    output n4436;
    output n4440;
    output n4442;
    output n4441;
    output n4444;
    output n4443;
    output n4446;
    output n4445;
    output [9:0]PWMdut_m4;
    output [9:0]PWMdut_m3;
    output [9:0]PWMdut_m2;
    output n4448;
    output n4447;
    output n4450;
    output n4449;
    output [9:0]PWMdut_m1;
    output n4452;
    output n4451;
    output n4454;
    output n4453;
    output n4456;
    output n4455;
    input \speed_avg_m4[3] ;
    output n4458;
    output n4457;
    output n4460;
    output n4459;
    output n4461;
    input \speed_avg_m4[12] ;
    input \speed_avg_m4[9] ;
    input \speed_avg_m4[8] ;
    output n4415;
    output n4414;
    
    wire clk_N_683 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    
    wire n22083, n21342;
    wire [28:0]backOut0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(77[9:17])
    wire [28:0]backOut1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(78[9:17])
    wire [28:0]n581;
    wire [20:0]subIn2_24__N_1340;
    wire [15:0]n1286;
    
    wire n30, n16394, clk_N_683_enable_392, n14334, n15696, n42, 
        n5304, n1061, n3832;
    wire [28:0]addOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(92[9:15])
    wire [28:0]intgOut0_28__N_1433;
    wire [28:0]intgOut0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(67[9:17])
    
    wire clk_N_683_enable_387, n14222, n21293, n21294, n7_c, n21295, 
        n5302, n21298, n21317, n21297, n56, n16270, n15694, n49;
    wire [21:0]n2581;
    
    wire clk_N_683_enable_70;
    wire [28:0]Out3_28__N_982;
    
    wire n16470, n8, n5300, clk_N_683_enable_42, n21377, n21344;
    wire [28:0]intgOut1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(68[9:17])
    wire [28:0]intgOut2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(69[9:17])
    wire [28:0]n641;
    
    wire n21296, n4328, n22084, n21383;
    wire [4:0]ss;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(96[9:11])
    wire [28:0]multOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(88[9:16])
    wire [53:0]multOut_28__N_1217;
    
    wire n5298, n18132;
    wire [21:0]n2341;
    
    wire n18133, n18360, n18361, n18359, n16260, n18029, n5400, 
        n5402, n18030, n35, n18028, n5396, n5398, n5296;
    wire [28:0]Out0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(72[9:13])
    
    wire clk_N_683_enable_98;
    wire [28:0]Out1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(73[9:13])
    
    wire clk_N_683_enable_126;
    wire [28:0]Out2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(74[9:13])
    
    wire clk_N_683_enable_154;
    wire [28:0]Out3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(75[9:13])
    
    wire clk_N_683_enable_182;
    wire [28:0]backOut2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(79[9:17])
    
    wire clk_N_683_enable_210;
    wire [28:0]backOut3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(80[9:17])
    
    wire clk_N_683_enable_238, n21321, n9;
    wire [28:0]n551;
    wire [24:0]subOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(84[9:15])
    
    wire n5767, n5769, n18358, n18357, n18583, n18584;
    wire [15:0]n1349;
    
    wire n18057, n5771, n5773, n18356, n18056;
    wire [15:0]n1328;
    
    wire n5775, n5777, n21341, n4, n3720, n16540, n5294, n18355, 
        n3624, n4_adj_2134, n16216, n4_adj_2135, n3768, n16544, 
        n4_adj_2136, n3672, n16536, n18354, n5292, n5779, n22105, 
        n21333, clk_N_683_enable_303, n14312, n5781, n5290, n5783, 
        clk_N_683_enable_331, n14284, n5785, n5787, n5789, n21334, 
        clk_N_683_enable_390, n14256, n5791, n21243, n21337, n18353, 
        n5793, n1, n18055, n14228, n5795, n21359, n14, n18352, 
        n18131, n4372, n4371, n19513, n18351, n18350, n5797, n5288, 
        n21382, n5799, n15, n19508, n11489, n5801, n5286, n5284, 
        n5803, n5807, n5480, n5282, n11439, n2533;
    wire [28:0]n671;
    
    wire n5278, n18027, n5392, n5394, n21299, n5350, n5318;
    wire [28:0]intgOut3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(70[9:17])
    
    wire n14307, n18130, n4374, n4373, n18054, n18129, n4376, 
        n4375, n5330, n5320, n5358, n5316, n5314, n5312, n5324, 
        n5310, n5308, n5362, n19420, n5306, n5356;
    wire [9:0]n2249;
    wire [9:0]n1399;
    
    wire n5354, n18349, n18128, n4378, n4377, n9_adj_2137, n9_adj_2138, 
        n5342, n18348, n18347, n18346, n21308, n22082;
    wire [20:0]n367;
    
    wire n5328, n18345, n3600, n21310, n5346, n19440, n5344, n21346;
    wire [20:0]subIn2_24__N_1156;
    
    wire n5340, n5334, n22099, n5332, n5280, n5338, n18053, n18344, 
        n5360, n5352, n16214;
    wire [28:0]backOut3_28__N_1678;
    
    wire n5348, n5326, n5336, n14_adj_2139, n10, n6, n18026, n5388, 
        n5390, n18025, n5384, n5386, n21353, n21311, n18024, n5380, 
        n5382, n18023, n5376, n5378, n18022, n5372, n5374, n18018, 
        n18019;
    wire [15:0]n1307;
    
    wire n30_adj_2140, n14343, n21312, n18020, n18021, n18017, n5370, 
        n21351;
    wire [9:0]n2261;
    wire [9:0]n1443;
    
    wire n21313, subIn1_24__N_1339, dirout_m3_N_1753, subIn1_24__N_1155, 
        dirout_m4_N_1756;
    wire [28:0]backOut2_28__N_1649;
    
    wire n18052;
    wire [28:0]Out2_28__N_953;
    wire [28:0]n121;
    wire [23:0]multIn2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(87[9:16])
    
    wire mult_29s_25s_0_pp_1_2, mult_29s_25s_0_pp_2_4, mult_29s_25s_0_pp_3_6, 
        mult_29s_25s_0_pp_4_8, mult_29s_25s_0_pp_5_10, mult_29s_25s_0_pp_6_12, 
        mult_29s_25s_0_pp_7_14, mult_29s_25s_0_pp_8_16, mult_29s_25s_0_pp_9_18, 
        mult_29s_25s_0_pp_10_20, mult_29s_25s_0_pp_11_22, mult_29s_25s_0_pp_12_24, 
        mult_29s_25s_0_pp_12_25, mult_29s_25s_0_pp_12_26, mult_29s_25s_0_pp_12_27, 
        mult_29s_25s_0_pp_12_28, mult_29s_25s_0_cin_lr_2, mult_29s_25s_0_cin_lr_4, 
        mult_29s_25s_0_cin_lr_6, mult_29s_25s_0_cin_lr_8, mult_29s_25s_0_cin_lr_10, 
        mult_29s_25s_0_cin_lr_12, mult_29s_25s_0_cin_lr_14, mult_29s_25s_0_cin_lr_16, 
        mult_29s_25s_0_cin_lr_18, mult_29s_25s_0_cin_lr_20, mult_29s_25s_0_cin_lr_22, 
        co_mult_29s_25s_0_0_1, mult_29s_25s_0_pp_0_2, co_mult_29s_25s_0_0_2, 
        s_mult_29s_25s_0_0_4, mult_29s_25s_0_pp_0_4, mult_29s_25s_0_pp_0_3, 
        mult_29s_25s_0_pp_1_4, mult_29s_25s_0_pp_1_3, co_mult_29s_25s_0_0_3, 
        s_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_6, mult_29s_25s_0_pp_0_6, 
        mult_29s_25s_0_pp_0_5, mult_29s_25s_0_pp_1_6, mult_29s_25s_0_pp_1_5, 
        co_mult_29s_25s_0_0_4, s_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_8, 
        mult_29s_25s_0_pp_0_8, mult_29s_25s_0_pp_0_7, mult_29s_25s_0_pp_1_8, 
        mult_29s_25s_0_pp_1_7, co_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_10, mult_29s_25s_0_pp_0_10, mult_29s_25s_0_pp_0_9, 
        mult_29s_25s_0_pp_1_10, mult_29s_25s_0_pp_1_9, co_mult_29s_25s_0_0_6, 
        s_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_12, mult_29s_25s_0_pp_0_12, 
        mult_29s_25s_0_pp_0_11, mult_29s_25s_0_pp_1_12, mult_29s_25s_0_pp_1_11, 
        co_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_14, 
        mult_29s_25s_0_pp_0_14, mult_29s_25s_0_pp_0_13, mult_29s_25s_0_pp_1_14, 
        mult_29s_25s_0_pp_1_13, co_mult_29s_25s_0_0_8, s_mult_29s_25s_0_0_15, 
        s_mult_29s_25s_0_0_16, mult_29s_25s_0_pp_0_16, mult_29s_25s_0_pp_0_15, 
        mult_29s_25s_0_pp_1_16, mult_29s_25s_0_pp_1_15, co_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_17, s_mult_29s_25s_0_0_18, mult_29s_25s_0_pp_0_18, 
        mult_29s_25s_0_pp_0_17, mult_29s_25s_0_pp_1_18, mult_29s_25s_0_pp_1_17, 
        co_mult_29s_25s_0_0_10, s_mult_29s_25s_0_0_19, s_mult_29s_25s_0_0_20, 
        mult_29s_25s_0_pp_0_20, mult_29s_25s_0_pp_0_19, mult_29s_25s_0_pp_1_20, 
        mult_29s_25s_0_pp_1_19, co_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_21, 
        s_mult_29s_25s_0_0_22, mult_29s_25s_0_pp_0_22, mult_29s_25s_0_pp_0_21, 
        mult_29s_25s_0_pp_1_22, mult_29s_25s_0_pp_1_21, co_mult_29s_25s_0_0_12, 
        s_mult_29s_25s_0_0_23, s_mult_29s_25s_0_0_24, mult_29s_25s_0_pp_0_24, 
        mult_29s_25s_0_pp_0_23, mult_29s_25s_0_pp_1_24, mult_29s_25s_0_pp_1_23, 
        co_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_25, s_mult_29s_25s_0_0_26, 
        mult_29s_25s_0_pp_0_26, mult_29s_25s_0_pp_0_25, mult_29s_25s_0_pp_1_26, 
        mult_29s_25s_0_pp_1_25, s_mult_29s_25s_0_0_27, s_mult_29s_25s_0_0_28, 
        mult_29s_25s_0_pp_0_28, mult_29s_25s_0_pp_0_27, mult_29s_25s_0_pp_1_28, 
        mult_29s_25s_0_pp_1_27, co_mult_29s_25s_0_1_1, s_mult_29s_25s_0_1_6, 
        mult_29s_25s_0_pp_2_6, co_mult_29s_25s_0_1_2, s_mult_29s_25s_0_1_7, 
        s_mult_29s_25s_0_1_8, mult_29s_25s_0_pp_2_8, mult_29s_25s_0_pp_2_7, 
        mult_29s_25s_0_pp_3_8, mult_29s_25s_0_pp_3_7, co_mult_29s_25s_0_1_3, 
        s_mult_29s_25s_0_1_9, s_mult_29s_25s_0_1_10, mult_29s_25s_0_pp_2_10, 
        mult_29s_25s_0_pp_2_9, mult_29s_25s_0_pp_3_10, mult_29s_25s_0_pp_3_9, 
        co_mult_29s_25s_0_1_4, s_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_12, 
        mult_29s_25s_0_pp_2_12, mult_29s_25s_0_pp_2_11, mult_29s_25s_0_pp_3_12, 
        mult_29s_25s_0_pp_3_11, co_mult_29s_25s_0_1_5, s_mult_29s_25s_0_1_13, 
        s_mult_29s_25s_0_1_14, mult_29s_25s_0_pp_2_14, mult_29s_25s_0_pp_2_13, 
        mult_29s_25s_0_pp_3_14, mult_29s_25s_0_pp_3_13, co_mult_29s_25s_0_1_6, 
        s_mult_29s_25s_0_1_15, s_mult_29s_25s_0_1_16, mult_29s_25s_0_pp_2_16, 
        mult_29s_25s_0_pp_2_15, mult_29s_25s_0_pp_3_16, mult_29s_25s_0_pp_3_15, 
        co_mult_29s_25s_0_1_7, s_mult_29s_25s_0_1_17, s_mult_29s_25s_0_1_18, 
        mult_29s_25s_0_pp_2_18, mult_29s_25s_0_pp_2_17, mult_29s_25s_0_pp_3_18, 
        mult_29s_25s_0_pp_3_17, co_mult_29s_25s_0_1_8, s_mult_29s_25s_0_1_19, 
        s_mult_29s_25s_0_1_20, mult_29s_25s_0_pp_2_20, mult_29s_25s_0_pp_2_19, 
        mult_29s_25s_0_pp_3_20, mult_29s_25s_0_pp_3_19, co_mult_29s_25s_0_1_9, 
        s_mult_29s_25s_0_1_21, s_mult_29s_25s_0_1_22, mult_29s_25s_0_pp_2_22, 
        mult_29s_25s_0_pp_2_21, mult_29s_25s_0_pp_3_22, mult_29s_25s_0_pp_3_21, 
        co_mult_29s_25s_0_1_10, s_mult_29s_25s_0_1_23, s_mult_29s_25s_0_1_24, 
        mult_29s_25s_0_pp_2_24, mult_29s_25s_0_pp_2_23, mult_29s_25s_0_pp_3_24, 
        mult_29s_25s_0_pp_3_23, co_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_25, 
        s_mult_29s_25s_0_1_26, mult_29s_25s_0_pp_2_26, mult_29s_25s_0_pp_2_25, 
        mult_29s_25s_0_pp_3_26, mult_29s_25s_0_pp_3_25, s_mult_29s_25s_0_1_27, 
        s_mult_29s_25s_0_1_28, mult_29s_25s_0_pp_2_28, mult_29s_25s_0_pp_2_27, 
        mult_29s_25s_0_pp_3_28, mult_29s_25s_0_pp_3_27, co_mult_29s_25s_0_2_1, 
        s_mult_29s_25s_0_2_10, mult_29s_25s_0_pp_4_10, co_mult_29s_25s_0_2_2, 
        s_mult_29s_25s_0_2_12, s_mult_29s_25s_0_2_11, mult_29s_25s_0_pp_4_12, 
        mult_29s_25s_0_pp_4_11, mult_29s_25s_0_pp_5_12, mult_29s_25s_0_pp_5_11, 
        co_mult_29s_25s_0_2_3, s_mult_29s_25s_0_2_13, s_mult_29s_25s_0_2_14, 
        mult_29s_25s_0_pp_4_14, mult_29s_25s_0_pp_4_13, mult_29s_25s_0_pp_5_14, 
        mult_29s_25s_0_pp_5_13, co_mult_29s_25s_0_2_4, s_mult_29s_25s_0_2_15, 
        s_mult_29s_25s_0_2_16, mult_29s_25s_0_pp_4_16, mult_29s_25s_0_pp_4_15, 
        mult_29s_25s_0_pp_5_16, mult_29s_25s_0_pp_5_15, co_mult_29s_25s_0_2_5, 
        s_mult_29s_25s_0_2_17, s_mult_29s_25s_0_2_18, mult_29s_25s_0_pp_4_18, 
        mult_29s_25s_0_pp_4_17, mult_29s_25s_0_pp_5_18, mult_29s_25s_0_pp_5_17, 
        co_mult_29s_25s_0_2_6, s_mult_29s_25s_0_2_19, s_mult_29s_25s_0_2_20, 
        mult_29s_25s_0_pp_4_20, mult_29s_25s_0_pp_4_19, mult_29s_25s_0_pp_5_20, 
        mult_29s_25s_0_pp_5_19, co_mult_29s_25s_0_2_7, s_mult_29s_25s_0_2_21, 
        s_mult_29s_25s_0_2_22, mult_29s_25s_0_pp_4_22, mult_29s_25s_0_pp_4_21, 
        mult_29s_25s_0_pp_5_22, mult_29s_25s_0_pp_5_21, co_mult_29s_25s_0_2_8, 
        s_mult_29s_25s_0_2_23, s_mult_29s_25s_0_2_24, mult_29s_25s_0_pp_4_24, 
        mult_29s_25s_0_pp_4_23, mult_29s_25s_0_pp_5_24, mult_29s_25s_0_pp_5_23, 
        co_mult_29s_25s_0_2_9, s_mult_29s_25s_0_2_25, s_mult_29s_25s_0_2_26, 
        mult_29s_25s_0_pp_4_26, mult_29s_25s_0_pp_4_25, mult_29s_25s_0_pp_5_26, 
        mult_29s_25s_0_pp_5_25, s_mult_29s_25s_0_2_27, s_mult_29s_25s_0_2_28, 
        mult_29s_25s_0_pp_4_28, mult_29s_25s_0_pp_4_27, mult_29s_25s_0_pp_5_28, 
        mult_29s_25s_0_pp_5_27, co_mult_29s_25s_0_3_1, s_mult_29s_25s_0_3_14, 
        mult_29s_25s_0_pp_6_14, co_mult_29s_25s_0_3_2, s_mult_29s_25s_0_3_15, 
        s_mult_29s_25s_0_3_16, mult_29s_25s_0_pp_6_16, mult_29s_25s_0_pp_6_15, 
        mult_29s_25s_0_pp_7_16, mult_29s_25s_0_pp_7_15, co_mult_29s_25s_0_3_3, 
        s_mult_29s_25s_0_3_17, s_mult_29s_25s_0_3_18, mult_29s_25s_0_pp_6_18, 
        mult_29s_25s_0_pp_6_17, mult_29s_25s_0_pp_7_18, mult_29s_25s_0_pp_7_17, 
        co_mult_29s_25s_0_3_4, s_mult_29s_25s_0_3_19, s_mult_29s_25s_0_3_20, 
        mult_29s_25s_0_pp_6_20, mult_29s_25s_0_pp_6_19, mult_29s_25s_0_pp_7_20, 
        mult_29s_25s_0_pp_7_19, co_mult_29s_25s_0_3_5, s_mult_29s_25s_0_3_21, 
        s_mult_29s_25s_0_3_22, mult_29s_25s_0_pp_6_22, mult_29s_25s_0_pp_6_21, 
        mult_29s_25s_0_pp_7_22, mult_29s_25s_0_pp_7_21, co_mult_29s_25s_0_3_6, 
        s_mult_29s_25s_0_3_23, s_mult_29s_25s_0_3_24, mult_29s_25s_0_pp_6_24, 
        mult_29s_25s_0_pp_6_23, mult_29s_25s_0_pp_7_24, mult_29s_25s_0_pp_7_23, 
        co_mult_29s_25s_0_3_7, s_mult_29s_25s_0_3_25, s_mult_29s_25s_0_3_26, 
        mult_29s_25s_0_pp_6_26, mult_29s_25s_0_pp_6_25, mult_29s_25s_0_pp_7_26, 
        mult_29s_25s_0_pp_7_25, s_mult_29s_25s_0_3_27, s_mult_29s_25s_0_3_28, 
        mult_29s_25s_0_pp_6_28, mult_29s_25s_0_pp_6_27, mult_29s_25s_0_pp_7_28, 
        mult_29s_25s_0_pp_7_27, co_mult_29s_25s_0_4_1, s_mult_29s_25s_0_4_18, 
        mult_29s_25s_0_pp_8_18, co_mult_29s_25s_0_4_2, s_mult_29s_25s_0_4_20, 
        s_mult_29s_25s_0_4_19, mult_29s_25s_0_pp_8_20, mult_29s_25s_0_pp_8_19, 
        mult_29s_25s_0_pp_9_20, mult_29s_25s_0_pp_9_19, co_mult_29s_25s_0_4_3, 
        s_mult_29s_25s_0_4_21, s_mult_29s_25s_0_4_22, mult_29s_25s_0_pp_8_22, 
        mult_29s_25s_0_pp_8_21, mult_29s_25s_0_pp_9_22, mult_29s_25s_0_pp_9_21, 
        co_mult_29s_25s_0_4_4, s_mult_29s_25s_0_4_23, s_mult_29s_25s_0_4_24, 
        mult_29s_25s_0_pp_8_24, mult_29s_25s_0_pp_8_23, mult_29s_25s_0_pp_9_24, 
        mult_29s_25s_0_pp_9_23, co_mult_29s_25s_0_4_5, s_mult_29s_25s_0_4_25, 
        s_mult_29s_25s_0_4_26, mult_29s_25s_0_pp_8_26, mult_29s_25s_0_pp_8_25, 
        mult_29s_25s_0_pp_9_26, mult_29s_25s_0_pp_9_25, s_mult_29s_25s_0_4_27, 
        s_mult_29s_25s_0_4_28, mult_29s_25s_0_pp_8_28, mult_29s_25s_0_pp_8_27, 
        mult_29s_25s_0_pp_9_28, mult_29s_25s_0_pp_9_27, co_mult_29s_25s_0_5_1, 
        s_mult_29s_25s_0_5_22, mult_29s_25s_0_pp_10_22, co_mult_29s_25s_0_5_2, 
        s_mult_29s_25s_0_5_23, s_mult_29s_25s_0_5_24, mult_29s_25s_0_pp_10_24, 
        mult_29s_25s_0_pp_10_23, mult_29s_25s_0_pp_11_24, mult_29s_25s_0_pp_11_23, 
        co_mult_29s_25s_0_5_3, s_mult_29s_25s_0_5_25, s_mult_29s_25s_0_5_26, 
        mult_29s_25s_0_pp_10_26, mult_29s_25s_0_pp_10_25, mult_29s_25s_0_pp_11_26, 
        mult_29s_25s_0_pp_11_25, s_mult_29s_25s_0_5_27, s_mult_29s_25s_0_5_28, 
        mult_29s_25s_0_pp_10_28, mult_29s_25s_0_pp_10_27, mult_29s_25s_0_pp_11_28, 
        mult_29s_25s_0_pp_11_27, co_mult_29s_25s_0_6_1, s_mult_29s_25s_0_6_24, 
        co_mult_29s_25s_0_6_2, s_mult_29s_25s_0_6_25, s_mult_29s_25s_0_6_26, 
        s_mult_29s_25s_0_6_27, s_mult_29s_25s_0_6_28, co_mult_29s_25s_0_7_1, 
        co_mult_29s_25s_0_7_2, mult_29s_25s_0_pp_2_5, co_mult_29s_25s_0_7_3, 
        s_mult_29s_25s_0_7_8, co_mult_29s_25s_0_7_4, s_mult_29s_25s_0_7_9, 
        s_mult_29s_25s_0_7_10, co_mult_29s_25s_0_7_5, s_mult_29s_25s_0_7_11, 
        s_mult_29s_25s_0_7_12, co_mult_29s_25s_0_7_6, s_mult_29s_25s_0_7_13, 
        s_mult_29s_25s_0_7_14, co_mult_29s_25s_0_7_7, s_mult_29s_25s_0_7_15, 
        s_mult_29s_25s_0_7_16, co_mult_29s_25s_0_7_8, s_mult_29s_25s_0_7_17, 
        s_mult_29s_25s_0_7_18, co_mult_29s_25s_0_7_9, s_mult_29s_25s_0_7_19, 
        s_mult_29s_25s_0_7_20, co_mult_29s_25s_0_7_10, s_mult_29s_25s_0_7_21, 
        s_mult_29s_25s_0_7_22, co_mult_29s_25s_0_7_11, s_mult_29s_25s_0_7_23, 
        s_mult_29s_25s_0_7_24, co_mult_29s_25s_0_7_12, s_mult_29s_25s_0_7_25, 
        s_mult_29s_25s_0_7_26, s_mult_29s_25s_0_7_27, s_mult_29s_25s_0_7_28, 
        co_mult_29s_25s_0_8_1, s_mult_29s_25s_0_8_12, co_mult_29s_25s_0_8_2, 
        s_mult_29s_25s_0_8_13, s_mult_29s_25s_0_8_14, mult_29s_25s_0_pp_6_13, 
        co_mult_29s_25s_0_8_3, s_mult_29s_25s_0_8_15, s_mult_29s_25s_0_8_16, 
        co_mult_29s_25s_0_8_4, s_mult_29s_25s_0_8_17, s_mult_29s_25s_0_8_18, 
        co_mult_29s_25s_0_8_5, s_mult_29s_25s_0_8_19, s_mult_29s_25s_0_8_20, 
        co_mult_29s_25s_0_8_6, s_mult_29s_25s_0_8_21, s_mult_29s_25s_0_8_22, 
        co_mult_29s_25s_0_8_7, s_mult_29s_25s_0_8_23, s_mult_29s_25s_0_8_24, 
        co_mult_29s_25s_0_8_8, s_mult_29s_25s_0_8_25, s_mult_29s_25s_0_8_26, 
        s_mult_29s_25s_0_8_27, s_mult_29s_25s_0_8_28, co_mult_29s_25s_0_9_1, 
        s_mult_29s_25s_0_9_20, co_mult_29s_25s_0_9_2, s_mult_29s_25s_0_9_21, 
        s_mult_29s_25s_0_9_22, mult_29s_25s_0_pp_10_21, co_mult_29s_25s_0_9_3, 
        s_mult_29s_25s_0_9_24, s_mult_29s_25s_0_9_23, co_mult_29s_25s_0_9_4, 
        s_mult_29s_25s_0_9_25, s_mult_29s_25s_0_9_26, s_mult_29s_25s_0_9_27, 
        s_mult_29s_25s_0_9_28, n30_adj_2141;
    wire [9:0]n2273;
    wire [9:0]n1487;
    
    wire co_mult_29s_25s_0_10_1, co_mult_29s_25s_0_10_2, mult_29s_25s_0_pp_4_9, 
        co_mult_29s_25s_0_10_3, co_mult_29s_25s_0_10_4, co_mult_29s_25s_0_10_5, 
        s_mult_29s_25s_0_10_16, co_mult_29s_25s_0_10_6, s_mult_29s_25s_0_10_17, 
        s_mult_29s_25s_0_10_18, co_mult_29s_25s_0_10_7, s_mult_29s_25s_0_10_19, 
        s_mult_29s_25s_0_10_20, co_mult_29s_25s_0_10_8, s_mult_29s_25s_0_10_21, 
        s_mult_29s_25s_0_10_22, co_mult_29s_25s_0_10_9, s_mult_29s_25s_0_10_23, 
        s_mult_29s_25s_0_10_24, co_mult_29s_25s_0_10_10, s_mult_29s_25s_0_10_25, 
        s_mult_29s_25s_0_10_26, s_mult_29s_25s_0_10_27, s_mult_29s_25s_0_10_28, 
        co_mult_29s_25s_0_11_1, s_mult_29s_25s_0_11_24, co_mult_29s_25s_0_11_2, 
        s_mult_29s_25s_0_11_25, s_mult_29s_25s_0_11_26, s_mult_29s_25s_0_11_27, 
        s_mult_29s_25s_0_11_28, co_t_mult_29s_25s_0_12_1, co_t_mult_29s_25s_0_12_2, 
        mult_29s_25s_0_pp_8_17, co_t_mult_29s_25s_0_12_3, co_t_mult_29s_25s_0_12_4, 
        co_t_mult_29s_25s_0_12_5, co_t_mult_29s_25s_0_12_6, mult_29s_25s_0_cin_lr_0, 
        mco, mco_1, mco_2, mco_3, mco_4, mco_5, mco_6, mco_7, 
        mco_8, mco_9, mco_10, mco_11, mco_12, mco_14, mco_15, 
        mco_16, mco_17, mco_18, mco_19, mco_20, mco_21, mco_22, 
        mco_23, mco_24, mco_25, mco_28, mco_29, mco_30, mco_31, 
        mco_32, mco_33, mco_34, mco_35, mco_36, mco_37, mco_38, 
        mco_42, mco_43, mco_44, mco_45, mco_46, mco_47, mco_48, 
        mco_49, mco_50, mco_51, mco_56, mco_57, mco_58, mco_59, 
        mco_60, mco_61, mco_62, mco_63, mco_64, mco_70, mco_71, 
        mco_72, mco_73, mco_74, mco_75, mco_76, mco_77, mco_84, 
        mco_85, mco_86, mco_87, mco_88, mco_89, mco_90, mco_98, 
        mco_99, mco_100, mco_101, mco_102, mco_103, mco_112, mco_113, 
        mco_114, mco_115, mco_116, mco_126, mco_127, mco_128, mco_129, 
        mco_140, mco_141, mco_142, mco_154, mco_155, n22093, n22094, 
        n35_adj_2142, n40, n36, n38, n32, n9_adj_2143, n7_adj_2144, 
        n30_adj_2145, n10_adj_2146, n8_adj_2147, n4_adj_2148, n9_adj_2149, 
        n7_adj_2150, n10_adj_2151, n8_adj_2152, n4_adj_2153, n9_adj_2154, 
        n7_adj_2155, n10_adj_2156, n8_adj_2157, n4_adj_2158, n9_adj_2159, 
        n7_adj_2160, n10_adj_2161, n8_adj_2162, n4_adj_2163, n14352, 
        n21356, n14338, n14_adj_2164, n10_adj_2165, n18568, n6_adj_2166, 
        n18569, n14_adj_2167, n10_adj_2168, n18505, n19534, n3648, 
        n35_adj_2169, n40_adj_2170, n36_adj_2171, n38_adj_2172, n32_adj_2173, 
        n18051, n34, n24, n18492, n18127, n4380, n4379, n3744, 
        n35_adj_2174, n40_adj_2175, n36_adj_2176, n6_adj_2177, n18506, 
        n18343, n18126, n4382, n4381, n38_adj_2178, n32_adj_2179, 
        n18125, n4384, n4383, n34_adj_2180, n24_adj_2181, n18124, 
        n4386, n4385, n14_adj_2182, n10_adj_2183, n18586, n18123, 
        n4388, n4387, n18050, n18342, n4389, n6_adj_2184, n18587, 
        n18049, n18048, n18047, n18046, n16212, n18341, n18045, 
        n18340, n3696, n35_adj_2185, n40_adj_2186, n36_adj_2187, n18044, 
        n38_adj_2188, n32_adj_2189, n18043, n34_adj_2190, n24_adj_2191, 
        n18339, n14361, n18338, n18337, n18336, n18042, n18041, 
        n18335, n18040, n18039, n18038, n18334, n18333, n18332, 
        n18331, n18037, n18036, n18330, n18329, n18328, n18253, 
        n18252, n18327, n18326, n18251, n18325, n18250, n18249, 
        n18035, n18248, n18034, n18033, n18324, n18323, n18247, 
        n18322, n18321, n18246, n18245, n18032, n5410, n14278, 
        n34_adj_2192, n24_adj_2193, n18320, n5408, n5406, n5404, 
        n18244, n18319, n18318, n5768, n5770, n5772, n5774, n5776, 
        n5778, n5780, n5782, n5784, n5786, n5788, n5790, n5792, 
        n5794, n5796, n5798, n5800, n5802, n5804, n5808, n5481;
    wire [28:0]n611;
    wire [28:0]addIn2_28__N_1375;
    
    wire n20045;
    wire [28:0]addIn2_28__N_1246;
    wire [9:0]n2285;
    wire [9:0]n1531;
    
    wire n18243, n20272, n18242, n18317, n20019, n18241, n18316, 
        n18315, n18240, n18314, n18239, n18238, n18313, n21378, 
        n18237, n21320, n18236, n18031, n18235, n18312, n14250, 
        n21379, n18311, n21325, n18234, n18310, n18149, n18233, 
        n18148, n18309, n18308, n18231, n16396, n18147, n18230, 
        n18434, n18433, n18432, n18431, n18430, n18429, n21326, 
        n18428, n18427, n18426, n18425, n18424, n18423, n18422, 
        n18421, n18420, n18419, n18418, n18417, n18416, n18415, 
        n18414, n18413, n18412, n18411, n18410, n18409, n18408, 
        n18407, n18406, n18405, n18404, n18403, n18402, n18401, 
        n18400, n18399, n18398, n18397, n18396, n18229, n18395, 
        n18146, n18145, n18394, n18228, n18393, n18227, n18392, 
        n18226, n18144, n20022, n18143, n18225, n21392, n18224, 
        n18391, n18390, n18389, n18142, n21391, n18223, n21388, 
        n18388, n21389, n21398, n21397, n18387, n18141, n18140, 
        n18386, n18385, n18222, n18221, n18220, n18139, n18219, 
        n18384, n18138, n18137, n18383, n18382, n18381, n18380, 
        n18379, n18378, n18377, n18376, n18375, n18374, n18373, 
        n18372, n18371, n18370, n18369, n18368, n18367, n18366, 
        n18365, n18364, n18064, n18063, n18062, n18061, n18136, 
        n18135, n18218, n18363, n18060, n18059, n18058, n18362;
    
    LUT4 mux_136_i11_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[10]), 
         .D(backOut1[10]), .Z(n581[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i6_4_lut (.A(\speed_avg_m4[5] ), .B(\speed_avg_m3[5] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i6_4_lut.init = 16'hcac0;
    LUT4 i11764_3_lut_4_lut (.A(n1286[15]), .B(n30), .C(n16394), .D(clk_N_683_enable_392), 
         .Z(n14334)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(346[7:42])
    defparam i11764_3_lut_4_lut.init = 16'hf700;
    LUT4 mux_136_i10_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[9]), 
         .D(backOut1[9]), .Z(n581[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i13_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[12]), 
         .D(speed_set_m3[12]), .Z(n5304)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_189_i19_3_lut_3_lut (.A(n1061), .B(n3832), .C(addOut[18]), 
         .Z(intgOut0_28__N_1433[18])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i19_3_lut_3_lut.init = 16'hbaba;
    FD1P3IX intgOut0_i0 (.D(addOut[0]), .SP(clk_N_683_enable_387), .CD(n14222), 
            .CK(clk_N_683), .Q(intgOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i0.GSR = "ENABLED";
    LUT4 i2_4_lut_4_lut (.A(n21293), .B(n21294), .C(n7_c), .D(n21295), 
         .Z(n18938)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam i2_4_lut_4_lut.init = 16'h4000;
    LUT4 mux_1186_i12_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[11]), 
         .D(speed_set_m3[11]), .Z(n5302)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i2_4_lut (.A(n21298), .B(n21317), .C(n21297), .D(n56), .Z(n16270)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'hfbfa;
    LUT4 mux_1241_i19_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[18]), 
         .D(speed_set_m4[18]), .Z(n2581[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i19_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i11_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[10]), 
         .D(speed_set_m4[10]), .Z(n2581[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_136_i8_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[7]), 
         .D(backOut1[7]), .Z(n581[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i6_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[5]), 
         .D(backOut1[5]), .Z(n581[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i4_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[3]), 
         .D(backOut1[3]), .Z(n581[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i4_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX backOut0_i0_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i0.GSR = "DISABLED";
    LUT4 mux_1241_i5_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[4]), 
         .D(speed_set_m4[4]), .Z(n2581[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i5_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3_2_lut_3_lut (.A(n21317), .B(n56), .C(n16470), .Z(n8)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i3_2_lut_3_lut.init = 16'he0e0;
    LUT4 mux_92_i19_4_lut (.A(\speed_avg_m4[18] ), .B(\speed_avg_m3[18] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i19_4_lut.init = 16'hcac0;
    LUT4 mux_136_i2_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[1]), 
         .D(backOut1[1]), .Z(n581[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i11_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[10]), 
         .D(speed_set_m3[10]), .Z(n5300)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i11_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX backOut1_i0_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i0.GSR = "DISABLED";
    LUT4 mux_136_i16_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[15]), 
         .D(backOut1[15]), .Z(n581[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_138_i21_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[20]), 
         .D(intgOut2[20]), .Z(n641[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i20_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[19]), 
         .D(intgOut2[19]), .Z(n641[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i20_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13672_2_lut_rep_315 (.A(n15696), .B(n42), .Z(n21296)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13672_2_lut_rep_315.init = 16'heeee;
    LUT4 mux_138_i19_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[18]), 
         .D(intgOut2[18]), .Z(n641[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i19_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i14_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[13]), 
         .D(intgOut2[13]), .Z(n641[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i14_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_92_i5_4_lut (.A(\speed_avg_m4[4] ), .B(\speed_avg_m3[4] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i5_4_lut.init = 16'hcac0;
    LUT4 mux_138_i13_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[12]), 
         .D(intgOut2[12]), .Z(n641[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_92_i4_3_lut (.A(\speed_avg_m3[3] ), .B(\speed_avg_m2[3] ), 
         .C(n4328), .Z(subIn2_24__N_1340[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i4_3_lut.init = 16'hcaca;
    LUT4 mux_138_i11_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[10]), 
         .D(intgOut2[10]), .Z(n641[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 i2_4_lut_adj_48 (.A(n22083), .B(n22084), .C(n21383), .D(ss[2]), 
         .Z(n4328)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i2_4_lut_adj_48.init = 16'h0322;
    LUT4 mux_92_i3_4_lut (.A(\speed_avg_m4[2] ), .B(\speed_avg_m3[2] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i3_4_lut.init = 16'hcac0;
    FD1S3AX multOut_i0 (.D(multOut_28__N_1217[0]), .CK(clk_N_683), .Q(multOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i0.GSR = "ENABLED";
    LUT4 mux_138_i5_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[4]), 
         .D(intgOut2[4]), .Z(n641[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i5_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i4_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[3]), 
         .D(intgOut2[3]), .Z(n641[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i23_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[22]), 
         .D(intgOut2[22]), .Z(n641[22])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i23_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1186_i10_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[9]), 
         .D(speed_set_m3[9]), .Z(n5298)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i1_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[0]), 
         .D(intgOut2[0]), .Z(n641[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_92_i2_4_lut (.A(\speed_avg_m4[1] ), .B(\speed_avg_m3[1] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i2_4_lut.init = 16'hcac0;
    LUT4 mux_138_i22_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[21]), 
         .D(intgOut2[21]), .Z(n641[21])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i22_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i17_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[16]), 
         .D(intgOut2[16]), .Z(n641[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i17_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i16_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[15]), 
         .D(intgOut2[15]), .Z(n641[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i9_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[8]), 
         .D(intgOut2[8]), .Z(n641[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i9_3_lut_4_lut.init = 16'hfe10;
    CCU2D sub_16_rep_3_add_2_21 (.A0(n2341[19]), .B0(n7), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18132), .COUT(n18133), .S0(n4417), .S1(n4416));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_21.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_21.INIT1 = 16'h5555;
    defparam sub_16_rep_3_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_21.INJECT1_1 = "NO";
    CCU2D add_15001_11 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18360), .COUT(n18361));
    defparam add_15001_11.INIT0 = 16'hf555;
    defparam add_15001_11.INIT1 = 16'hf555;
    defparam add_15001_11.INJECT1_0 = "NO";
    defparam add_15001_11.INJECT1_1 = "NO";
    LUT4 mux_138_i6_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[5]), 
         .D(intgOut2[5]), .Z(n641[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i6_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15001_9 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18359), .COUT(n18360));
    defparam add_15001_9.INIT0 = 16'hf555;
    defparam add_15001_9.INIT1 = 16'h0aaa;
    defparam add_15001_9.INJECT1_0 = "NO";
    defparam add_15001_9.INJECT1_1 = "NO";
    LUT4 mux_138_i3_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[2]), 
         .D(intgOut2[2]), .Z(n641[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i2_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[1]), 
         .D(intgOut2[1]), .Z(n641[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i2_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13708_2_lut_3_lut_4_lut (.A(n15696), .B(n42), .C(n49), .D(n15694), 
         .Z(n16260)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i13708_2_lut_3_lut_4_lut.init = 16'heee0;
    LUT4 mux_92_i1_4_lut (.A(\speed_avg_m4[0] ), .B(\speed_avg_m3[0] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i1_4_lut.init = 16'hcac0;
    LUT4 mux_136_i13_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[12]), 
         .D(backOut1[12]), .Z(n581[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_138_i8_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[7]), 
         .D(intgOut2[7]), .Z(n641[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i8_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1176_17 (.A0(n5400), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5402), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18029), 
          .COUT(n18030), .S0(n2341[15]), .S1(n2341[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_17.INIT0 = 16'hf555;
    defparam add_1176_17.INIT1 = 16'hf555;
    defparam add_1176_17.INJECT1_0 = "NO";
    defparam add_1176_17.INJECT1_1 = "NO";
    LUT4 mux_138_i12_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[11]), 
         .D(intgOut2[11]), .Z(n641[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i12_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i24_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[23]), 
         .D(intgOut2[23]), .Z(n641[23])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i24_3_lut_4_lut.init = 16'hfe10;
    LUT4 i17112_2_lut_rep_312_2_lut_3_lut_4_lut (.A(n16470), .B(n35), .C(n42), 
         .D(n15696), .Z(n21293)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))))) */ ;
    defparam i17112_2_lut_rep_312_2_lut_3_lut_4_lut.init = 16'h111f;
    CCU2D add_1176_15 (.A0(n5396), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5398), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18028), 
          .COUT(n18029), .S0(n2341[13]), .S1(n2341[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_15.INIT0 = 16'hf555;
    defparam add_1176_15.INIT1 = 16'hf555;
    defparam add_1176_15.INJECT1_0 = "NO";
    defparam add_1176_15.INJECT1_1 = "NO";
    LUT4 mux_136_i15_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[14]), 
         .D(backOut1[14]), .Z(n581[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_138_i25_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[24]), 
         .D(intgOut2[24]), .Z(n641[24])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1186_i9_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[8]), 
         .D(speed_set_m3[8]), .Z(n5296)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_138_i26_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[25]), 
         .D(intgOut2[25]), .Z(n641[25])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i26_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX Out0_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_98), .CK(clk_N_683), 
            .Q(Out0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i0.GSR = "ENABLED";
    FD1P3AX Out1_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_126), .CK(clk_N_683), 
            .Q(Out1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i0.GSR = "ENABLED";
    FD1P3AX Out2_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_154), .CK(clk_N_683), 
            .Q(Out2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i0.GSR = "ENABLED";
    FD1P3AX Out3_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_182), .CK(clk_N_683), 
            .Q(Out3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i0.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i0.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i0 (.D(Out3_28__N_982[0]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i0.GSR = "DISABLED";
    LUT4 mux_138_i7_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[6]), 
         .D(intgOut2[6]), .Z(n641[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_92_i18_4_lut (.A(\speed_avg_m4[17] ), .B(\speed_avg_m3[17] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i18_4_lut.init = 16'hcac0;
    LUT4 mux_135_i2_4_lut (.A(backOut2[1]), .B(backOut3[1]), .C(n21321), 
         .D(n9), .Z(n551[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i2_4_lut.init = 16'h0aca;
    LUT4 mux_138_i10_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[9]), 
         .D(intgOut2[9]), .Z(n641[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i10_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i15_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[14]), 
         .D(intgOut2[14]), .Z(n641[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i18_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[17]), 
         .D(intgOut2[17]), .Z(n641[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i18_3_lut_4_lut.init = 16'hfe10;
    FD1S3AX subOut_i0 (.D(\subOut_24__N_1177[0] ), .CK(clk_N_683), .Q(subOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i0.GSR = "ENABLED";
    LUT4 mux_138_i27_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[26]), 
         .D(intgOut2[26]), .Z(n641[26])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i27_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3285_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m2[1]), .Z(n5767)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3285_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i28_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[27]), 
         .D(intgOut2[27]), .Z(n641[27])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i28_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i29_3_lut_4_lut (.A(n21377), .B(n21344), .C(intgOut1[28]), 
         .D(intgOut2[28]), .Z(n641[28])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i29_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3287_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m2[2]), .Z(n5769)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3287_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15001_7 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18358), .COUT(n18359));
    defparam add_15001_7.INIT0 = 16'h0aaa;
    defparam add_15001_7.INIT1 = 16'hf555;
    defparam add_15001_7.INJECT1_0 = "NO";
    defparam add_15001_7.INJECT1_1 = "NO";
    CCU2D add_15001_5 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18357), .COUT(n18358));
    defparam add_15001_5.INIT0 = 16'h0aaa;
    defparam add_15001_5.INIT1 = 16'h0aaa;
    defparam add_15001_5.INJECT1_0 = "NO";
    defparam add_15001_5.INJECT1_1 = "NO";
    CCU2D add_223_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[13]), .B1(n18583), .C1(n18584), .D1(Out3[28]), .COUT(n18057), 
          .S1(n1349[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_1.INIT0 = 16'hF000;
    defparam add_223_1.INIT1 = 16'h56aa;
    defparam add_223_1.INJECT1_0 = "NO";
    defparam add_223_1.INJECT1_1 = "NO";
    LUT4 mux_136_i17_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[16]), 
         .D(backOut1[16]), .Z(n581[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3289_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m2[3]), .Z(n5771)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3289_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3291_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m2[4]), .Z(n5773)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3291_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15001_3 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18356), .COUT(n18357));
    defparam add_15001_3.INIT0 = 16'hf555;
    defparam add_15001_3.INIT1 = 16'hf555;
    defparam add_15001_3.INJECT1_0 = "NO";
    defparam add_15001_3.INJECT1_1 = "NO";
    LUT4 mux_136_i18_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[17]), 
         .D(backOut1[17]), .Z(n581[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i18_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_219_17 (.A0(Out2[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18056), 
          .S0(n1328[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_17.INIT0 = 16'h5aaa;
    defparam add_219_17.INIT1 = 16'h0000;
    defparam add_219_17.INJECT1_0 = "NO";
    defparam add_219_17.INJECT1_1 = "NO";
    LUT4 i3293_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m2[5]), .Z(n5775)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3293_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3295_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m2[6]), .Z(n5777)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3295_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_92_i17_4_lut (.A(\speed_avg_m4[16] ), .B(\speed_avg_m3[16] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i17_4_lut.init = 16'hcac0;
    CCU2D add_15001_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[4]), .B1(speed_set_m2[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18356));
    defparam add_15001_1.INIT0 = 16'hF000;
    defparam add_15001_1.INIT1 = 16'ha666;
    defparam add_15001_1.INJECT1_0 = "NO";
    defparam add_15001_1.INJECT1_1 = "NO";
    LUT4 i13975_3_lut_4_lut (.A(n21377), .B(n21341), .C(n4), .D(n3720), 
         .Z(n16540)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13975_3_lut_4_lut.init = 16'hfeee;
    LUT4 mux_1186_i8_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[7]), 
         .D(speed_set_m3[7]), .Z(n5294)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i8_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_15002_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18355), 
          .S0(n3624));
    defparam add_15002_cout.INIT0 = 16'h0000;
    defparam add_15002_cout.INIT1 = 16'h0000;
    defparam add_15002_cout.INJECT1_0 = "NO";
    defparam add_15002_cout.INJECT1_1 = "NO";
    LUT4 i13666_3_lut_4_lut (.A(n21377), .B(n21341), .C(n4_adj_2134), 
         .D(n3624), .Z(n16216)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13666_3_lut_4_lut.init = 16'hfeee;
    LUT4 mux_135_i3_4_lut (.A(backOut2[2]), .B(backOut3[2]), .C(n21321), 
         .D(n9), .Z(n551[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i3_4_lut.init = 16'h0aca;
    LUT4 mux_92_i16_4_lut (.A(\speed_avg_m4[15] ), .B(\speed_avg_m3[15] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i16_4_lut.init = 16'hcac0;
    LUT4 i13979_3_lut_4_lut (.A(n21377), .B(n21341), .C(n4_adj_2135), 
         .D(n3768), .Z(n16544)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13979_3_lut_4_lut.init = 16'hfeee;
    LUT4 mux_136_i19_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[18]), 
         .D(backOut1[18]), .Z(n581[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13971_3_lut_4_lut (.A(n21377), .B(n21341), .C(n4_adj_2136), 
         .D(n3672), .Z(n16536)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13971_3_lut_4_lut.init = 16'hfeee;
    LUT4 mux_92_i15_4_lut (.A(\speed_avg_m4[14] ), .B(\speed_avg_m3[14] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i15_4_lut.init = 16'hcac0;
    CCU2D add_15002_20 (.A0(speed_set_m1[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18354), .COUT(n18355));
    defparam add_15002_20.INIT0 = 16'h5aaa;
    defparam add_15002_20.INIT1 = 16'h0aaa;
    defparam add_15002_20.INJECT1_0 = "NO";
    defparam add_15002_20.INJECT1_1 = "NO";
    LUT4 mux_92_i14_4_lut (.A(\speed_avg_m4[13] ), .B(\speed_avg_m3[13] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i14_4_lut.init = 16'hcac0;
    LUT4 mux_136_i20_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[19]), 
         .D(backOut1[19]), .Z(n581[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i7_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[6]), 
         .D(speed_set_m3[6]), .Z(n5292)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i4_4_lut (.A(backOut2[3]), .B(backOut3[3]), .C(n21321), 
         .D(n9), .Z(n551[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i4_4_lut.init = 16'h0aca;
    LUT4 mux_136_i21_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[20]), 
         .D(backOut1[20]), .Z(n581[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3297_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m2[7]), .Z(n5779)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3297_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_136_i22_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[21]), 
         .D(backOut1[21]), .Z(n581[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11760_2_lut_3_lut_4_lut (.A(n22105), .B(n21333), .C(clk_N_683_enable_303), 
         .D(ss[1]), .Z(n14312)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11760_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i3299_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m2[8]), .Z(n5781)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3299_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1186_i6_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[5]), 
         .D(speed_set_m3[5]), .Z(n5290)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3301_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m2[9]), .Z(n5783)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3301_3_lut_4_lut.init = 16'hfe10;
    LUT4 i11732_2_lut_3_lut_4_lut (.A(n22105), .B(n21333), .C(clk_N_683_enable_331), 
         .D(ss[1]), .Z(n14284)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11732_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i3303_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m2[10]), .Z(n5785)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3303_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i5_4_lut (.A(backOut2[4]), .B(backOut3[4]), .C(n21321), 
         .D(n9), .Z(n551[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i5_4_lut.init = 16'h0aca;
    LUT4 i3305_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m2[11]), .Z(n5787)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3305_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_136_i23_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[22]), 
         .D(backOut1[22]), .Z(n581[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3307_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m2[12]), .Z(n5789)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3307_3_lut_4_lut.init = 16'hfe10;
    LUT4 i11704_2_lut_3_lut_4_lut (.A(n22105), .B(n21334), .C(clk_N_683_enable_390), 
         .D(ss[1]), .Z(n14256)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11704_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i3309_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m2[13]), .Z(n5791)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3309_3_lut_4_lut.init = 16'hfe10;
    PFUMX i17299 (.BLUT(n21243), .ALUT(n21337), .C0(n22105), .Z(clk_N_683_enable_154));
    CCU2D add_15002_18 (.A0(speed_set_m1[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18353), .COUT(n18354));
    defparam add_15002_18.INIT0 = 16'h5aaa;
    defparam add_15002_18.INIT1 = 16'h5aaa;
    defparam add_15002_18.INJECT1_0 = "NO";
    defparam add_15002_18.INJECT1_1 = "NO";
    LUT4 mux_136_i24_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[23]), 
         .D(backOut1[23]), .Z(n581[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3311_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m2[14]), .Z(n5793)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3311_3_lut_4_lut.init = 16'hfe10;
    FD1S3IX ss_i0 (.D(n1), .CK(clk_N_683), .CD(ss[4]), .Q(ss[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i0.GSR = "ENABLED";
    CCU2D add_219_15 (.A0(Out2[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18055), 
          .COUT(n18056), .S0(n1328[13]), .S1(n1328[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_15.INIT0 = 16'h5aaa;
    defparam add_219_15.INIT1 = 16'h5aaa;
    defparam add_219_15.INJECT1_0 = "NO";
    defparam add_219_15.INJECT1_1 = "NO";
    LUT4 i11676_2_lut_3_lut_4_lut (.A(n22105), .B(n21334), .C(clk_N_683_enable_387), 
         .D(ss[1]), .Z(n14228)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11676_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i3313_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m2[15]), .Z(n5795)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3313_3_lut_4_lut.init = 16'hfe10;
    FD1S3IX ss_i1 (.D(n21359), .CK(clk_N_683), .CD(ss[4]), .Q(ss[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i1.GSR = "ENABLED";
    FD1S3IX ss_i2 (.D(n14), .CK(clk_N_683), .CD(ss[4]), .Q(ss[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i2.GSR = "ENABLED";
    CCU2D add_15002_16 (.A0(speed_set_m1[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18352), .COUT(n18353));
    defparam add_15002_16.INIT0 = 16'h5aaa;
    defparam add_15002_16.INIT1 = 16'h5aaa;
    defparam add_15002_16.INJECT1_0 = "NO";
    defparam add_15002_16.INJECT1_1 = "NO";
    LUT4 mux_136_i25_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[24]), 
         .D(backOut1[24]), .Z(n581[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i25_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_16_rep_3_add_2_19 (.A0(n2341[17]), .B0(n4372), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[18]), .B1(n4371), .C1(GND_net), .D1(GND_net), 
          .CIN(n18131), .COUT(n18132), .S0(n4419), .S1(n4418));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_19.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_19.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_19.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(n21337), .B(n22105), .C(n19513), .D(ss[3]), 
         .Z(clk_N_683_enable_126)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam i1_4_lut_4_lut.init = 16'hb888;
    CCU2D add_15002_14 (.A0(speed_set_m1[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18351), .COUT(n18352));
    defparam add_15002_14.INIT0 = 16'h5555;
    defparam add_15002_14.INIT1 = 16'h5aaa;
    defparam add_15002_14.INJECT1_0 = "NO";
    defparam add_15002_14.INJECT1_1 = "NO";
    CCU2D add_15002_12 (.A0(speed_set_m1[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18350), .COUT(n18351));
    defparam add_15002_12.INIT0 = 16'h5aaa;
    defparam add_15002_12.INIT1 = 16'h5aaa;
    defparam add_15002_12.INJECT1_0 = "NO";
    defparam add_15002_12.INJECT1_1 = "NO";
    LUT4 i3315_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m2[16]), .Z(n5797)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3315_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_136_i26_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[25]), 
         .D(backOut1[25]), .Z(n581[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i5_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[4]), 
         .D(speed_set_m3[4]), .Z(n5288)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i6_4_lut (.A(backOut2[5]), .B(backOut3[5]), .C(n21321), 
         .D(n9), .Z(n551[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i6_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_4_lut_adj_49 (.A(n21337), .B(n22105), .C(n21382), .D(n21383), 
         .Z(clk_N_683_enable_98)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B+((D)+!C))) */ ;
    defparam i1_4_lut_4_lut_adj_49.init = 16'h88b8;
    LUT4 i3317_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m2[17]), .Z(n5799)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3317_3_lut_4_lut.init = 16'hfe10;
    FD1S3IX ss_i3 (.D(n15), .CK(clk_N_683), .CD(ss[4]), .Q(ss[3]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i3.GSR = "ENABLED";
    LUT4 mux_92_i13_3_lut (.A(\speed_avg_m3[12] ), .B(\speed_avg_m2[12] ), 
         .C(n4328), .Z(subIn2_24__N_1340[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i13_3_lut.init = 16'hcaca;
    LUT4 mux_136_i27_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[26]), 
         .D(backOut1[26]), .Z(n581[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut (.A(n21337), .B(n22105), .C(n22100), .Z(n19508)) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i1_4_lut_4_lut_adj_50 (.A(n21337), .B(n22105), .C(n11489), .D(ss[3]), 
         .Z(clk_N_683_enable_182)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B+!(C (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_50.init = 16'hb888;
    LUT4 i3319_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m2[18]), .Z(n5801)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3319_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_136_i28_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[27]), 
         .D(backOut1[27]), .Z(n581[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i4_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[3]), 
         .D(speed_set_m3[3]), .Z(n5286)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1186_i3_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[2]), 
         .D(speed_set_m3[2]), .Z(n5284)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3321_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m2[19]), .Z(n5803)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3321_3_lut_4_lut.init = 16'hfe10;
    LUT4 i3325_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m2[20]), .Z(n5807)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i3325_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_135_i7_4_lut (.A(backOut2[6]), .B(backOut3[6]), .C(n21321), 
         .D(n9), .Z(n551[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i7_4_lut.init = 16'h0aca;
    LUT4 mux_136_i29_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[28]), 
         .D(backOut1[28]), .Z(n581[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2998_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m2[0]), .Z(n5480)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam i2998_3_lut_4_lut.init = 16'hfe10;
    LUT4 i52_2_lut_rep_316 (.A(n15694), .B(n49), .Z(n21297)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(138[23] 139[51])
    defparam i52_2_lut_rep_316.init = 16'h4444;
    LUT4 mux_136_i1_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[0]), 
         .D(backOut1[0]), .Z(n581[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i2_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[1]), 
         .D(speed_set_m3[1]), .Z(n5282)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n15694), .B(n49), .C(n11439), .D(n21298), 
         .Z(n2533)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(138[23] 139[51])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf040;
    LUT4 i1_2_lut_rep_317 (.A(n15696), .B(n42), .Z(n21298)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam i1_2_lut_rep_317.init = 16'h4444;
    LUT4 mux_135_i8_4_lut (.A(backOut2[7]), .B(backOut3[7]), .C(n21321), 
         .D(n9), .Z(n551[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i8_4_lut.init = 16'h0aca;
    LUT4 mux_139_i27_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[26]), 
         .D(n641[26]), .Z(n671[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i1_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[0]), 
         .D(speed_set_m3[0]), .Z(n5278)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i1_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_1176_13 (.A0(n5392), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5394), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18027), 
          .COUT(n18028), .S0(n2341[11]), .S1(n2341[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_13.INIT0 = 16'hf555;
    defparam add_1176_13.INIT1 = 16'hf555;
    defparam add_1176_13.INJECT1_0 = "NO";
    defparam add_1176_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_318 (.A(n16470), .B(n35), .Z(n21299)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam i1_2_lut_rep_318.init = 16'h4444;
    LUT4 mux_92_i12_4_lut (.A(\speed_avg_m4[11] ), .B(\speed_avg_m3[11] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i12_4_lut.init = 16'hcac0;
    LUT4 mux_135_i9_4_lut (.A(backOut2[8]), .B(backOut3[8]), .C(n21321), 
         .D(n9), .Z(n551[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i9_4_lut.init = 16'h0aca;
    LUT4 mux_92_i11_4_lut (.A(\speed_avg_m4[10] ), .B(\speed_avg_m3[10] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i11_4_lut.init = 16'hcac0;
    LUT4 mux_139_i22_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[21]), 
         .D(n641[21]), .Z(n671[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i21_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[20]), 
         .D(n641[20]), .Z(n671[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i20_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[19]), 
         .D(n641[19]), .Z(n671[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i18_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[17]), 
         .D(n641[17]), .Z(n671[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1185_i15_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m4[14]), .Z(n5350)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i10_4_lut (.A(backOut2[9]), .B(backOut3[9]), .C(n21321), 
         .D(n9), .Z(n551[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i10_4_lut.init = 16'h0aca;
    LUT4 mux_139_i16_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[15]), 
         .D(n641[15]), .Z(n671[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i14_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[13]), 
         .D(n641[13]), .Z(n671[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i20_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[19]), 
         .D(speed_set_m3[19]), .Z(n5318)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_92_i10_3_lut (.A(\speed_avg_m3[9] ), .B(\speed_avg_m2[9] ), 
         .C(n4328), .Z(subIn2_24__N_1340[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i10_3_lut.init = 16'hcaca;
    FD1P3IX intgOut3_i0 (.D(addOut[0]), .SP(clk_N_683_enable_303), .CD(n14307), 
            .CK(clk_N_683), .Q(intgOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i0.GSR = "ENABLED";
    CCU2D sub_16_rep_3_add_2_17 (.A0(n2341[15]), .B0(n4374), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[16]), .B1(n4373), .C1(GND_net), .D1(GND_net), 
          .CIN(n18130), .COUT(n18131), .S0(n4421), .S1(n4420));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_17.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_17.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_17.INJECT1_1 = "NO";
    LUT4 mux_92_i9_3_lut (.A(\speed_avg_m3[8] ), .B(\speed_avg_m2[8] ), 
         .C(n4328), .Z(subIn2_24__N_1340[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i9_3_lut.init = 16'hcaca;
    LUT4 mux_136_i9_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[8]), 
         .D(backOut1[8]), .Z(n581[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i9_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_219_13 (.A0(Out2[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18054), 
          .COUT(n18055), .S0(n1328[11]), .S1(n1328[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_13.INIT0 = 16'h5aaa;
    defparam add_219_13.INIT1 = 16'h5aaa;
    defparam add_219_13.INJECT1_0 = "NO";
    defparam add_219_13.INJECT1_1 = "NO";
    LUT4 mux_139_i13_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[12]), 
         .D(n641[12]), .Z(n671[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i13_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_16_rep_3_add_2_15 (.A0(n2341[13]), .B0(n4376), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[14]), .B1(n4375), .C1(GND_net), .D1(GND_net), 
          .CIN(n18129), .COUT(n18130), .S0(n4423), .S1(n4422));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_15.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_15.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_15.INJECT1_1 = "NO";
    LUT4 mux_136_i7_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[6]), 
         .D(backOut1[6]), .Z(n581[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i10_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[9]), 
         .D(n641[9]), .Z(n671[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i7_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[6]), 
         .D(n641[6]), .Z(n671[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1185_i5_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m4[4]), .Z(n5330)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i11_4_lut (.A(backOut2[10]), .B(backOut3[10]), .C(n21321), 
         .D(n9), .Z(n551[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i11_4_lut.init = 16'h0aca;
    LUT4 mux_139_i6_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[5]), 
         .D(n641[5]), .Z(n671[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i5_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[4]), 
         .D(n641[4]), .Z(n671[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i26_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[25]), 
         .D(n641[25]), .Z(n671[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i21_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[20]), 
         .D(speed_set_m3[20]), .Z(n5320)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i19_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m4[18]), .Z(n5358)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1186_i19_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[18]), 
         .D(speed_set_m3[18]), .Z(n5316)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1186_i18_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[17]), 
         .D(speed_set_m3[17]), .Z(n5314)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_139_i24_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[23]), 
         .D(n641[23]), .Z(n671[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i12_4_lut (.A(backOut2[11]), .B(backOut3[11]), .C(n21321), 
         .D(n9), .Z(n551[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i12_4_lut.init = 16'h0aca;
    LUT4 mux_1186_i17_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[16]), 
         .D(speed_set_m3[16]), .Z(n5312)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_139_i23_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[22]), 
         .D(n641[22]), .Z(n671[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i1_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[0]), 
         .D(n641[0]), .Z(n671[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i5_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[4]), 
         .D(backOut1[4]), .Z(n581[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1185_i2_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m4[1]), .Z(n5324)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_136_i3_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[2]), 
         .D(backOut1[2]), .Z(n581[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i19_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[18]), 
         .D(n641[18]), .Z(n671[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i17_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[16]), 
         .D(n641[16]), .Z(n671[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1186_i16_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[15]), 
         .D(speed_set_m3[15]), .Z(n5310)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1186_i15_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[14]), 
         .D(speed_set_m3[14]), .Z(n5308)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_139_i15_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[14]), 
         .D(n641[14]), .Z(n671[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1185_i21_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m4[20]), .Z(n5362)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_139_i12_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[11]), 
         .D(n641[11]), .Z(n671[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i11_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[10]), 
         .D(n641[10]), .Z(n671[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i8_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[7]), 
         .D(n641[7]), .Z(n671[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i8_3_lut_4_lut.init = 16'hfd20;
    FD1S3AY ss_i4_rep_414 (.D(n19420), .CK(clk_N_683), .Q(n22105));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i4_rep_414.GSR = "ENABLED";
    LUT4 mux_1186_i14_3_lut_4_lut (.A(n15696), .B(n42), .C(speed_set_m2[13]), 
         .D(speed_set_m3[13]), .Z(n5306)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1186_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_136_i14_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[13]), 
         .D(backOut1[13]), .Z(n581[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i8_3_lut (.A(\speed_avg_m3[7] ), .B(\speed_avg_m2[7] ), 
         .C(n4328), .Z(subIn2_24__N_1340[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i8_3_lut.init = 16'hcaca;
    LUT4 mux_139_i3_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[2]), 
         .D(n641[2]), .Z(n671[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1185_i18_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m4[17]), .Z(n5356)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_136_i12_3_lut_4_lut (.A(n22083), .B(n21342), .C(backOut0[11]), 
         .D(backOut1[11]), .Z(n581[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i9_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[8]), 
         .D(n641[8]), .Z(n671[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_135_i13_4_lut (.A(backOut2[12]), .B(backOut3[12]), .C(n21321), 
         .D(n9), .Z(n551[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i13_4_lut.init = 16'h0aca;
    LUT4 mux_139_i2_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[1]), 
         .D(n641[1]), .Z(n671[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i7_4_lut (.A(\speed_avg_m4[6] ), .B(\speed_avg_m3[6] ), 
         .C(n21328), .D(n4322), .Z(subIn2_24__N_1340[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i7_4_lut.init = 16'hcac0;
    LUT4 mux_139_i25_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[24]), 
         .D(n641[24]), .Z(n671[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_230_i4_3_lut_4_lut_3_lut (.A(n30), .B(n1286[15]), .C(n2249[3]), 
         .Z(n1399[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(346[25:42])
    defparam mux_230_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_139_i4_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[3]), 
         .D(n641[3]), .Z(n671[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1185_i17_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m4[16]), .Z(n5354)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i17_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_15002_10 (.A0(speed_set_m1[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18349), .COUT(n18350));
    defparam add_15002_10.INIT0 = 16'h5555;
    defparam add_15002_10.INIT1 = 16'h5555;
    defparam add_15002_10.INJECT1_0 = "NO";
    defparam add_15002_10.INJECT1_1 = "NO";
    LUT4 mux_139_i28_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[27]), 
         .D(n641[27]), .Z(n671[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i28_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_16_rep_3_add_2_13 (.A0(n2341[11]), .B0(n4378), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[12]), .B1(n4377), .C1(GND_net), .D1(GND_net), 
          .CIN(n18128), .COUT(n18129), .S0(n4425), .S1(n4424));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_13.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_13.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_13.INJECT1_1 = "NO";
    LUT4 mux_139_i29_3_lut_4_lut (.A(n22083), .B(n21341), .C(intgOut0[28]), 
         .D(n641[28]), .Z(n671[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2_3_lut_rep_336_4_lut (.A(n22083), .B(n21344), .C(n9_adj_2137), 
         .D(n9_adj_2138), .Z(n21317)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(170[9:16])
    defparam i2_3_lut_rep_336_4_lut.init = 16'hd000;
    LUT4 mux_1185_i11_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m4[10]), .Z(n5342)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i11_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_15002_8 (.A0(speed_set_m1[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18348), .COUT(n18349));
    defparam add_15002_8.INIT0 = 16'h5aaa;
    defparam add_15002_8.INIT1 = 16'h5555;
    defparam add_15002_8.INJECT1_0 = "NO";
    defparam add_15002_8.INJECT1_1 = "NO";
    CCU2D add_15002_6 (.A0(speed_set_m1[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18347), .COUT(n18348));
    defparam add_15002_6.INIT0 = 16'h5aaa;
    defparam add_15002_6.INIT1 = 16'h5aaa;
    defparam add_15002_6.INJECT1_0 = "NO";
    defparam add_15002_6.INJECT1_1 = "NO";
    CCU2D add_15002_4 (.A0(speed_set_m1[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18346), .COUT(n18347));
    defparam add_15002_4.INIT0 = 16'h5555;
    defparam add_15002_4.INIT1 = 16'h5aaa;
    defparam add_15002_4.INJECT1_0 = "NO";
    defparam add_15002_4.INJECT1_1 = "NO";
    CCU2D add_15002_2 (.A0(speed_set_m1[1]), .B0(speed_set_m1[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18346));
    defparam add_15002_2.INIT0 = 16'h1000;
    defparam add_15002_2.INIT1 = 16'h5555;
    defparam add_15002_2.INJECT1_0 = "NO";
    defparam add_15002_2.INJECT1_1 = "NO";
    LUT4 mux_91_i8_3_lut_4_lut_4_lut (.A(n21308), .B(\speed_avg_m4[7] ), 
         .C(n4322), .D(n22082), .Z(n367[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i8_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_1185_i4_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m4[3]), .Z(n5328)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i14_4_lut (.A(backOut2[13]), .B(backOut3[13]), .C(n21321), 
         .D(n9), .Z(n551[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i14_4_lut.init = 16'h0aca;
    CCU2D add_15003_17 (.A0(speed_set_m1[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18345), .S1(n3600));
    defparam add_15003_17.INIT0 = 16'h5555;
    defparam add_15003_17.INIT1 = 16'h0000;
    defparam add_15003_17.INJECT1_0 = "NO";
    defparam add_15003_17.INJECT1_1 = "NO";
    LUT4 mux_230_i9_3_lut_4_lut_3_lut (.A(n30), .B(n1286[15]), .C(n2249[8]), 
         .Z(n1399[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(346[25:42])
    defparam mux_230_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i11653_3_lut_4_lut (.A(n1061), .B(n3832), .C(n21310), .D(clk_N_683_enable_387), 
         .Z(n14222)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i11653_3_lut_4_lut.init = 16'hfe00;
    LUT4 mux_1185_i13_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m4[12]), .Z(n5346)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i15_4_lut (.A(backOut2[14]), .B(backOut3[14]), .C(n21321), 
         .D(n9), .Z(n551[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i15_4_lut.init = 16'h0aca;
    LUT4 mux_230_i6_3_lut_4_lut_3_lut (.A(n30), .B(n1286[15]), .C(n2249[5]), 
         .Z(n1399[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(346[25:42])
    defparam mux_230_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i1_4_lut (.A(ss[1]), .B(n19508), .C(n22105), .D(n19440), .Z(clk_N_683_enable_210)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hc4c0;
    LUT4 mux_1185_i12_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m4[11]), .Z(n5344)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i2_3_lut (.A(ss[3]), .B(ss[2]), .C(ss[0]), .Z(n19440)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_3_lut.init = 16'h2020;
    LUT4 subIn2_24__I_25_i19_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[18] ), 
         .D(\speed_avg_m2[18] ), .Z(subIn2_24__N_1156[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i10_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m4[9]), .Z(n5340)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i7_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m4[6]), .Z(n5334)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i16_4_lut (.A(backOut2[15]), .B(backOut3[15]), .C(n21321), 
         .D(n9), .Z(n551[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i16_4_lut.init = 16'h0aca;
    FD1S3IX ss_i2_rep_408 (.D(n14), .CK(clk_N_683), .CD(ss[4]), .Q(n22099));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i2_rep_408.GSR = "ENABLED";
    LUT4 subIn2_24__I_25_i18_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[17] ), 
         .D(\speed_avg_m2[17] ), .Z(subIn2_24__N_1156[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i17_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[16] ), 
         .D(\speed_avg_m2[16] ), .Z(subIn2_24__N_1156[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i16_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[15] ), 
         .D(\speed_avg_m2[15] ), .Z(subIn2_24__N_1156[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13141_2_lut_rep_402 (.A(ss[1]), .B(ss[0]), .Z(n21383)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13141_2_lut_rep_402.init = 16'heeee;
    LUT4 subIn2_24__I_25_i15_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[14] ), 
         .D(\speed_avg_m2[14] ), .Z(subIn2_24__N_1156[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i6_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m4[5]), .Z(n5332)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13834_2_lut_3_lut_4_lut (.A(ss[1]), .B(ss[0]), .C(ss[3]), .D(n22099), 
         .Z(n16394)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13834_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_51 (.A(ss[1]), .B(n19508), .C(n22105), .D(n19440), 
         .Z(clk_N_683_enable_238)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_51.init = 16'hc8c0;
    LUT4 subIn2_24__I_25_i14_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[13] ), 
         .D(\speed_avg_m2[13] ), .Z(subIn2_24__N_1156[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i13_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[12] ), 
         .D(subIn2_24__N_1340[12]), .Z(subIn2_24__N_1156[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i1_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m4[0]), .Z(n5280)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i12_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[11] ), 
         .D(\speed_avg_m2[11] ), .Z(subIn2_24__N_1156[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i11_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[10] ), 
         .D(\speed_avg_m2[10] ), .Z(subIn2_24__N_1156[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i10_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[9] ), 
         .D(subIn2_24__N_1340[9]), .Z(subIn2_24__N_1156[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i9_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[8] ), 
         .D(subIn2_24__N_1340[8]), .Z(subIn2_24__N_1156[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_230_i10_3_lut_4_lut_3_lut (.A(n30), .B(n1286[15]), .C(n2249[9]), 
         .Z(n1399[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(346[25:42])
    defparam mux_230_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_230_i7_3_lut_4_lut_3_lut (.A(n30), .B(n1286[15]), .C(n2249[6]), 
         .Z(n1399[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(346[25:42])
    defparam mux_230_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 subIn2_24__I_25_i8_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[7] ), 
         .D(subIn2_24__N_1340[7]), .Z(subIn2_24__N_1156[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i9_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m4[8]), .Z(n5338)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i9_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_219_11 (.A0(Out2[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18053), 
          .COUT(n18054), .S0(n1328[9]), .S1(n1328[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_11.INIT0 = 16'h5aaa;
    defparam add_219_11.INIT1 = 16'h5aaa;
    defparam add_219_11.INJECT1_0 = "NO";
    defparam add_219_11.INJECT1_1 = "NO";
    CCU2D add_15003_15 (.A0(speed_set_m1[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18344), .COUT(n18345));
    defparam add_15003_15.INIT0 = 16'hf555;
    defparam add_15003_15.INIT1 = 16'hf555;
    defparam add_15003_15.INJECT1_0 = "NO";
    defparam add_15003_15.INJECT1_1 = "NO";
    LUT4 mux_135_i17_4_lut (.A(backOut2[16]), .B(backOut3[16]), .C(n21321), 
         .D(n9), .Z(n551[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i17_4_lut.init = 16'h0aca;
    LUT4 subIn2_24__I_25_i7_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[6] ), 
         .D(\speed_avg_m2[6] ), .Z(subIn2_24__N_1156[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i20_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m4[19]), .Z(n5360)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i6_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[5] ), 
         .D(\speed_avg_m2[5] ), .Z(subIn2_24__N_1156[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i16_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m4[15]), .Z(n5352)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_adj_52 (.A(n16216), .B(n16214), .C(n21337), .D(n22105), 
         .Z(clk_N_683_enable_387)) /* synthesis lut_function=((B (C (D))+!B (C+!(D)))+!A) */ ;
    defparam i1_4_lut_adj_52.init = 16'hf577;
    LUT4 i13368_2_lut (.A(addOut[16]), .B(n22105), .Z(backOut3_28__N_1678[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13368_2_lut.init = 16'h2222;
    LUT4 subIn2_24__I_25_i5_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[4] ), 
         .D(\speed_avg_m2[4] ), .Z(subIn2_24__N_1156[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i4_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[3] ), 
         .D(subIn2_24__N_1340[3]), .Z(subIn2_24__N_1156[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i3_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[2] ), 
         .D(\speed_avg_m2[2] ), .Z(subIn2_24__N_1156[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i2_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[1] ), 
         .D(\speed_avg_m2[1] ), .Z(subIn2_24__N_1156[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13068_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[19] ), 
         .D(\speed_avg_m2[19] ), .Z(n5)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i13068_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i1_3_lut_4_lut (.A(ss[2]), .B(n21346), .C(\speed_avg_m1[0] ), 
         .D(\speed_avg_m2[0] ), .Z(subIn2_24__N_1156[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i14_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m4[13]), .Z(n5348)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1185_i3_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m4[2]), .Z(n5326)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_135_i18_4_lut (.A(backOut2[17]), .B(backOut3[17]), .C(n21321), 
         .D(n9), .Z(n551[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i18_4_lut.init = 16'h0aca;
    LUT4 mux_1185_i8_3_lut_4_lut (.A(n16470), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m4[7]), .Z(n5336)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1185_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 i7_4_lut (.A(Out3[3]), .B(n14_adj_2139), .C(n10), .D(Out3[4]), 
         .Z(n18583)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut (.A(Out3[11]), .B(Out3[7]), .C(Out3[2]), .D(Out3[10]), 
         .Z(n14_adj_2139)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(Out3[9]), .B(Out3[1]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i4_4_lut (.A(Out3[5]), .B(Out3[6]), .C(Out3[0]), .D(n6), .Z(n18584)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(Out3[8]), .B(Out3[12]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i1_2_lut.init = 16'heeee;
    CCU2D add_1176_11 (.A0(n5388), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5390), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18026), 
          .COUT(n18027), .S0(n2341[9]), .S1(n2341[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_11.INIT0 = 16'hf555;
    defparam add_1176_11.INIT1 = 16'hf555;
    defparam add_1176_11.INJECT1_0 = "NO";
    defparam add_1176_11.INJECT1_1 = "NO";
    LUT4 mux_230_i8_3_lut_4_lut_3_lut (.A(n30), .B(n1286[15]), .C(n2249[7]), 
         .Z(n1399[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(346[25:42])
    defparam mux_230_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_135_i19_4_lut (.A(backOut2[18]), .B(backOut3[18]), .C(n21321), 
         .D(n9), .Z(n551[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i19_4_lut.init = 16'h0aca;
    CCU2D add_1176_9 (.A0(n5384), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5386), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18025), 
          .COUT(n18026), .S0(n2341[7]), .S1(n2341[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_9.INIT0 = 16'hf555;
    defparam add_1176_9.INIT1 = 16'hf555;
    defparam add_1176_9.INJECT1_0 = "NO";
    defparam add_1176_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_330_3_lut_4_lut (.A(ss[3]), .B(n21353), .C(ss[1]), 
         .D(n22105), .Z(n21311)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_330_3_lut_4_lut.init = 16'hfffd;
    CCU2D add_1176_7 (.A0(n5380), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5382), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18024), 
          .COUT(n18025), .S0(n2341[5]), .S1(n2341[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_7.INIT0 = 16'hf555;
    defparam add_1176_7.INIT1 = 16'hf555;
    defparam add_1176_7.INJECT1_0 = "NO";
    defparam add_1176_7.INJECT1_1 = "NO";
    CCU2D add_1176_5 (.A0(n5376), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5378), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18023), 
          .COUT(n18024), .S0(n2341[3]), .S1(n2341[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_5.INIT0 = 16'hf555;
    defparam add_1176_5.INIT1 = 16'hf555;
    defparam add_1176_5.INJECT1_0 = "NO";
    defparam add_1176_5.INJECT1_1 = "NO";
    CCU2D add_1176_3 (.A0(n5372), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5374), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18022), 
          .COUT(n18023), .S0(n2341[1]), .S1(n2341[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_3.INIT0 = 16'hf555;
    defparam add_1176_3.INIT1 = 16'hf555;
    defparam add_1176_3.INJECT1_0 = "NO";
    defparam add_1176_3.INJECT1_1 = "NO";
    CCU2D add_1170_5 (.A0(n1286[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1286[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18018), 
          .COUT(n18019), .S0(n2249[3]), .S1(n2249[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1170_5.INIT0 = 16'hf555;
    defparam add_1170_5.INIT1 = 16'hf555;
    defparam add_1170_5.INJECT1_0 = "NO";
    defparam add_1170_5.INJECT1_1 = "NO";
    LUT4 mux_135_i20_4_lut (.A(backOut2[19]), .B(backOut3[19]), .C(n21321), 
         .D(n9), .Z(n551[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i20_4_lut.init = 16'h0aca;
    LUT4 i11773_3_lut_4_lut (.A(n1307[15]), .B(n30_adj_2140), .C(n16394), 
         .D(clk_N_683_enable_392), .Z(n14343)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[7:42])
    defparam i11773_3_lut_4_lut.init = 16'hf700;
    LUT4 i1_2_lut_rep_331_3_lut_4_lut (.A(ss[3]), .B(n21353), .C(ss[1]), 
         .D(n22105), .Z(n21312)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_331_3_lut_4_lut.init = 16'hffdf;
    CCU2D add_1170_9 (.A0(n1286[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1286[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18020), 
          .COUT(n18021), .S0(n2249[7]), .S1(n2249[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1170_9.INIT0 = 16'hf555;
    defparam add_1170_9.INIT1 = 16'hf555;
    defparam add_1170_9.INJECT1_0 = "NO";
    defparam add_1170_9.INJECT1_1 = "NO";
    CCU2D add_1170_3 (.A0(n1286[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1286[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18017), 
          .COUT(n18018), .S0(n2249[1]), .S1(n2249[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1170_3.INIT0 = 16'hf555;
    defparam add_1170_3.INIT1 = 16'hf555;
    defparam add_1170_3.INJECT1_0 = "NO";
    defparam add_1170_3.INJECT1_1 = "NO";
    CCU2D add_1176_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5370), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18022), 
          .S1(n2341[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_1.INIT0 = 16'hF000;
    defparam add_1176_1.INIT1 = 16'h0aaa;
    defparam add_1176_1.INJECT1_0 = "NO";
    defparam add_1176_1.INJECT1_1 = "NO";
    CCU2D add_1170_7 (.A0(n1286[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1286[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18019), 
          .COUT(n18020), .S0(n2249[5]), .S1(n2249[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1170_7.INIT0 = 16'hf555;
    defparam add_1170_7.INIT1 = 16'hf555;
    defparam add_1170_7.INJECT1_0 = "NO";
    defparam add_1170_7.INJECT1_1 = "NO";
    CCU2D add_1170_11 (.A0(n1286[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18021), 
          .S0(n2249[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1170_11.INIT0 = 16'hf555;
    defparam add_1170_11.INIT1 = 16'h0000;
    defparam add_1170_11.INJECT1_0 = "NO";
    defparam add_1170_11.INJECT1_1 = "NO";
    CCU2D add_1170_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1286[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18017), 
          .S1(n2249[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1170_1.INIT0 = 16'hF000;
    defparam add_1170_1.INIT1 = 16'h0aaa;
    defparam add_1170_1.INJECT1_0 = "NO";
    defparam add_1170_1.INJECT1_1 = "NO";
    FD1S3AY ss_i4 (.D(n19420), .CK(clk_N_683), .Q(ss[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i4.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_329_3_lut_4_lut (.A(ss[2]), .B(n21351), .C(ss[1]), 
         .D(n22105), .Z(n21310)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_329_3_lut_4_lut.init = 16'hfffd;
    LUT4 mux_237_i4_3_lut_4_lut_3_lut (.A(n30_adj_2140), .B(n1307[15]), 
         .C(n2261[3]), .Z(n1443[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[25:42])
    defparam mux_237_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_135_i21_4_lut (.A(backOut2[20]), .B(backOut3[20]), .C(n21321), 
         .D(n9), .Z(n551[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i21_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_rep_332_3_lut_4_lut (.A(ss[2]), .B(n21351), .C(ss[1]), 
         .D(n22105), .Z(n21313)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_332_3_lut_4_lut.init = 16'hffdf;
    FD1P3AX dirout_m2_347 (.D(subIn1_24__N_1339), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m2_347.GSR = "DISABLED";
    FD1P3AX dirout_m3_348 (.D(dirout_m3_N_1753), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m3_348.GSR = "DISABLED";
    FD1P3AX dirout_m1_346 (.D(subIn1_24__N_1155), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m1_346.GSR = "DISABLED";
    FD1P3AX dirout_m4_349 (.D(dirout_m4_N_1756), .SP(clk_N_683_enable_392), 
            .CK(clk_N_683), .Q(dir_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m4_349.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i28.GSR = "DISABLED";
    CCU2D add_219_9 (.A0(Out2[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18052), 
          .COUT(n18053), .S0(n1328[7]), .S1(n1328[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_9.INIT0 = 16'h5aaa;
    defparam add_219_9.INIT1 = 16'h5aaa;
    defparam add_219_9.INJECT1_0 = "NO";
    defparam add_219_9.INJECT1_1 = "NO";
    FD1P3AX backOut1_i0_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_42), 
            .CK(clk_N_683), .Q(backOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i1.GSR = "DISABLED";
    LUT4 mux_237_i9_3_lut_4_lut_3_lut (.A(n30_adj_2140), .B(n1307[15]), 
         .C(n2261[8]), .Z(n1443[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[25:42])
    defparam mux_237_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FD1S3AX addOut_2081__i0 (.D(n121[0]), .CK(clk_N_683), .Q(addOut[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i0.GSR = "ENABLED";
    AND2 AND2_t64 (.A(subOut[0]), .B(GND_net), .Z(multOut_28__N_1217[0])) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1256[10:66])
    AND2 AND2_t61 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1262[10:66])
    AND2 AND2_t58 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1268[10:66])
    AND2 AND2_t55 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1274[10:66])
    AND2 AND2_t52 (.A(subOut[0]), .B(multIn2[4]), .Z(mult_29s_25s_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1280[10:66])
    AND2 AND2_t49 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_5_10)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1286[10:68])
    AND2 AND2_t46 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_6_12)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1292[10:68])
    AND2 AND2_t43 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_7_14)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1298[10:68])
    AND2 AND2_t40 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_8_16)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1304[10:68])
    AND2 AND2_t37 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_9_18)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1310[10:68])
    AND2 AND2_t34 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_10_20)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1316[10:69])
    AND2 AND2_t31 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_11_22)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1322[10:69])
    ND2 ND2_t28 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t27 (.A(subOut[1]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_25)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t26 (.A(subOut[2]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t25 (.A(subOut[3]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_27)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t24 (.A(subOut[4]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_12 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_14 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_16 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_18 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_20 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_22 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_0_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_0_2), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_1_2), .CI(GND_net), .COUT(co_mult_29s_25s_0_0_1), 
           .S1(multOut_28__N_1217[2])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_2 (.A0(mult_29s_25s_0_pp_0_3), .A1(mult_29s_25s_0_pp_0_4), 
           .B0(mult_29s_25s_0_pp_1_3), .B1(mult_29s_25s_0_pp_1_4), .CI(co_mult_29s_25s_0_0_1), 
           .COUT(co_mult_29s_25s_0_0_2), .S0(multOut_28__N_1217[3]), .S1(s_mult_29s_25s_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_3 (.A0(mult_29s_25s_0_pp_0_5), .A1(mult_29s_25s_0_pp_0_6), 
           .B0(mult_29s_25s_0_pp_1_5), .B1(mult_29s_25s_0_pp_1_6), .CI(co_mult_29s_25s_0_0_2), 
           .COUT(co_mult_29s_25s_0_0_3), .S0(s_mult_29s_25s_0_0_5), .S1(s_mult_29s_25s_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_4 (.A0(mult_29s_25s_0_pp_0_7), .A1(mult_29s_25s_0_pp_0_8), 
           .B0(mult_29s_25s_0_pp_1_7), .B1(mult_29s_25s_0_pp_1_8), .CI(co_mult_29s_25s_0_0_3), 
           .COUT(co_mult_29s_25s_0_0_4), .S0(s_mult_29s_25s_0_0_7), .S1(s_mult_29s_25s_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_5 (.A0(mult_29s_25s_0_pp_0_9), .A1(mult_29s_25s_0_pp_0_10), 
           .B0(mult_29s_25s_0_pp_1_9), .B1(mult_29s_25s_0_pp_1_10), .CI(co_mult_29s_25s_0_0_4), 
           .COUT(co_mult_29s_25s_0_0_5), .S0(s_mult_29s_25s_0_0_9), .S1(s_mult_29s_25s_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_6 (.A0(mult_29s_25s_0_pp_0_11), .A1(mult_29s_25s_0_pp_0_12), 
           .B0(mult_29s_25s_0_pp_1_11), .B1(mult_29s_25s_0_pp_1_12), .CI(co_mult_29s_25s_0_0_5), 
           .COUT(co_mult_29s_25s_0_0_6), .S0(s_mult_29s_25s_0_0_11), .S1(s_mult_29s_25s_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_7 (.A0(mult_29s_25s_0_pp_0_13), .A1(mult_29s_25s_0_pp_0_14), 
           .B0(mult_29s_25s_0_pp_1_13), .B1(mult_29s_25s_0_pp_1_14), .CI(co_mult_29s_25s_0_0_6), 
           .COUT(co_mult_29s_25s_0_0_7), .S0(s_mult_29s_25s_0_0_13), .S1(s_mult_29s_25s_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_8 (.A0(mult_29s_25s_0_pp_0_15), .A1(mult_29s_25s_0_pp_0_16), 
           .B0(mult_29s_25s_0_pp_1_15), .B1(mult_29s_25s_0_pp_1_16), .CI(co_mult_29s_25s_0_0_7), 
           .COUT(co_mult_29s_25s_0_0_8), .S0(s_mult_29s_25s_0_0_15), .S1(s_mult_29s_25s_0_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_9 (.A0(mult_29s_25s_0_pp_0_17), .A1(mult_29s_25s_0_pp_0_18), 
           .B0(mult_29s_25s_0_pp_1_17), .B1(mult_29s_25s_0_pp_1_18), .CI(co_mult_29s_25s_0_0_8), 
           .COUT(co_mult_29s_25s_0_0_9), .S0(s_mult_29s_25s_0_0_17), .S1(s_mult_29s_25s_0_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_10 (.A0(mult_29s_25s_0_pp_0_19), .A1(mult_29s_25s_0_pp_0_20), 
           .B0(mult_29s_25s_0_pp_1_19), .B1(mult_29s_25s_0_pp_1_20), .CI(co_mult_29s_25s_0_0_9), 
           .COUT(co_mult_29s_25s_0_0_10), .S0(s_mult_29s_25s_0_0_19), .S1(s_mult_29s_25s_0_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_11 (.A0(mult_29s_25s_0_pp_0_21), .A1(mult_29s_25s_0_pp_0_22), 
           .B0(mult_29s_25s_0_pp_1_21), .B1(mult_29s_25s_0_pp_1_22), .CI(co_mult_29s_25s_0_0_10), 
           .COUT(co_mult_29s_25s_0_0_11), .S0(s_mult_29s_25s_0_0_21), .S1(s_mult_29s_25s_0_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_12 (.A0(mult_29s_25s_0_pp_0_23), .A1(mult_29s_25s_0_pp_0_24), 
           .B0(mult_29s_25s_0_pp_1_23), .B1(mult_29s_25s_0_pp_1_24), .CI(co_mult_29s_25s_0_0_11), 
           .COUT(co_mult_29s_25s_0_0_12), .S0(s_mult_29s_25s_0_0_23), .S1(s_mult_29s_25s_0_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_13 (.A0(mult_29s_25s_0_pp_0_25), .A1(mult_29s_25s_0_pp_0_26), 
           .B0(mult_29s_25s_0_pp_1_25), .B1(mult_29s_25s_0_pp_1_26), .CI(co_mult_29s_25s_0_0_12), 
           .COUT(co_mult_29s_25s_0_0_13), .S0(s_mult_29s_25s_0_0_25), .S1(s_mult_29s_25s_0_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_14 (.A0(mult_29s_25s_0_pp_0_27), .A1(mult_29s_25s_0_pp_0_28), 
           .B0(mult_29s_25s_0_pp_1_27), .B1(mult_29s_25s_0_pp_1_28), .CI(co_mult_29s_25s_0_0_13), 
           .S0(s_mult_29s_25s_0_0_27), .S1(s_mult_29s_25s_0_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_1_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_2_6), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_3_6), .CI(GND_net), .COUT(co_mult_29s_25s_0_1_1), 
           .S1(s_mult_29s_25s_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_2 (.A0(mult_29s_25s_0_pp_2_7), .A1(mult_29s_25s_0_pp_2_8), 
           .B0(mult_29s_25s_0_pp_3_7), .B1(mult_29s_25s_0_pp_3_8), .CI(co_mult_29s_25s_0_1_1), 
           .COUT(co_mult_29s_25s_0_1_2), .S0(s_mult_29s_25s_0_1_7), .S1(s_mult_29s_25s_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_3 (.A0(mult_29s_25s_0_pp_2_9), .A1(mult_29s_25s_0_pp_2_10), 
           .B0(mult_29s_25s_0_pp_3_9), .B1(mult_29s_25s_0_pp_3_10), .CI(co_mult_29s_25s_0_1_2), 
           .COUT(co_mult_29s_25s_0_1_3), .S0(s_mult_29s_25s_0_1_9), .S1(s_mult_29s_25s_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_4 (.A0(mult_29s_25s_0_pp_2_11), .A1(mult_29s_25s_0_pp_2_12), 
           .B0(mult_29s_25s_0_pp_3_11), .B1(mult_29s_25s_0_pp_3_12), .CI(co_mult_29s_25s_0_1_3), 
           .COUT(co_mult_29s_25s_0_1_4), .S0(s_mult_29s_25s_0_1_11), .S1(s_mult_29s_25s_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_5 (.A0(mult_29s_25s_0_pp_2_13), .A1(mult_29s_25s_0_pp_2_14), 
           .B0(mult_29s_25s_0_pp_3_13), .B1(mult_29s_25s_0_pp_3_14), .CI(co_mult_29s_25s_0_1_4), 
           .COUT(co_mult_29s_25s_0_1_5), .S0(s_mult_29s_25s_0_1_13), .S1(s_mult_29s_25s_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_6 (.A0(mult_29s_25s_0_pp_2_15), .A1(mult_29s_25s_0_pp_2_16), 
           .B0(mult_29s_25s_0_pp_3_15), .B1(mult_29s_25s_0_pp_3_16), .CI(co_mult_29s_25s_0_1_5), 
           .COUT(co_mult_29s_25s_0_1_6), .S0(s_mult_29s_25s_0_1_15), .S1(s_mult_29s_25s_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_7 (.A0(mult_29s_25s_0_pp_2_17), .A1(mult_29s_25s_0_pp_2_18), 
           .B0(mult_29s_25s_0_pp_3_17), .B1(mult_29s_25s_0_pp_3_18), .CI(co_mult_29s_25s_0_1_6), 
           .COUT(co_mult_29s_25s_0_1_7), .S0(s_mult_29s_25s_0_1_17), .S1(s_mult_29s_25s_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_8 (.A0(mult_29s_25s_0_pp_2_19), .A1(mult_29s_25s_0_pp_2_20), 
           .B0(mult_29s_25s_0_pp_3_19), .B1(mult_29s_25s_0_pp_3_20), .CI(co_mult_29s_25s_0_1_7), 
           .COUT(co_mult_29s_25s_0_1_8), .S0(s_mult_29s_25s_0_1_19), .S1(s_mult_29s_25s_0_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_9 (.A0(mult_29s_25s_0_pp_2_21), .A1(mult_29s_25s_0_pp_2_22), 
           .B0(mult_29s_25s_0_pp_3_21), .B1(mult_29s_25s_0_pp_3_22), .CI(co_mult_29s_25s_0_1_8), 
           .COUT(co_mult_29s_25s_0_1_9), .S0(s_mult_29s_25s_0_1_21), .S1(s_mult_29s_25s_0_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_10 (.A0(mult_29s_25s_0_pp_2_23), .A1(mult_29s_25s_0_pp_2_24), 
           .B0(mult_29s_25s_0_pp_3_23), .B1(mult_29s_25s_0_pp_3_24), .CI(co_mult_29s_25s_0_1_9), 
           .COUT(co_mult_29s_25s_0_1_10), .S0(s_mult_29s_25s_0_1_23), .S1(s_mult_29s_25s_0_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_11 (.A0(mult_29s_25s_0_pp_2_25), .A1(mult_29s_25s_0_pp_2_26), 
           .B0(mult_29s_25s_0_pp_3_25), .B1(mult_29s_25s_0_pp_3_26), .CI(co_mult_29s_25s_0_1_10), 
           .COUT(co_mult_29s_25s_0_1_11), .S0(s_mult_29s_25s_0_1_25), .S1(s_mult_29s_25s_0_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_12 (.A0(mult_29s_25s_0_pp_2_27), .A1(mult_29s_25s_0_pp_2_28), 
           .B0(mult_29s_25s_0_pp_3_27), .B1(mult_29s_25s_0_pp_3_28), .CI(co_mult_29s_25s_0_1_11), 
           .S0(s_mult_29s_25s_0_1_27), .S1(s_mult_29s_25s_0_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_2_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_4_10), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_5_10), .CI(GND_net), .COUT(co_mult_29s_25s_0_2_1), 
           .S1(s_mult_29s_25s_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_2 (.A0(mult_29s_25s_0_pp_4_11), .A1(mult_29s_25s_0_pp_4_12), 
           .B0(mult_29s_25s_0_pp_5_11), .B1(mult_29s_25s_0_pp_5_12), .CI(co_mult_29s_25s_0_2_1), 
           .COUT(co_mult_29s_25s_0_2_2), .S0(s_mult_29s_25s_0_2_11), .S1(s_mult_29s_25s_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_3 (.A0(mult_29s_25s_0_pp_4_13), .A1(mult_29s_25s_0_pp_4_14), 
           .B0(mult_29s_25s_0_pp_5_13), .B1(mult_29s_25s_0_pp_5_14), .CI(co_mult_29s_25s_0_2_2), 
           .COUT(co_mult_29s_25s_0_2_3), .S0(s_mult_29s_25s_0_2_13), .S1(s_mult_29s_25s_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_4 (.A0(mult_29s_25s_0_pp_4_15), .A1(mult_29s_25s_0_pp_4_16), 
           .B0(mult_29s_25s_0_pp_5_15), .B1(mult_29s_25s_0_pp_5_16), .CI(co_mult_29s_25s_0_2_3), 
           .COUT(co_mult_29s_25s_0_2_4), .S0(s_mult_29s_25s_0_2_15), .S1(s_mult_29s_25s_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_5 (.A0(mult_29s_25s_0_pp_4_17), .A1(mult_29s_25s_0_pp_4_18), 
           .B0(mult_29s_25s_0_pp_5_17), .B1(mult_29s_25s_0_pp_5_18), .CI(co_mult_29s_25s_0_2_4), 
           .COUT(co_mult_29s_25s_0_2_5), .S0(s_mult_29s_25s_0_2_17), .S1(s_mult_29s_25s_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_6 (.A0(mult_29s_25s_0_pp_4_19), .A1(mult_29s_25s_0_pp_4_20), 
           .B0(mult_29s_25s_0_pp_5_19), .B1(mult_29s_25s_0_pp_5_20), .CI(co_mult_29s_25s_0_2_5), 
           .COUT(co_mult_29s_25s_0_2_6), .S0(s_mult_29s_25s_0_2_19), .S1(s_mult_29s_25s_0_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_7 (.A0(mult_29s_25s_0_pp_4_21), .A1(mult_29s_25s_0_pp_4_22), 
           .B0(mult_29s_25s_0_pp_5_21), .B1(mult_29s_25s_0_pp_5_22), .CI(co_mult_29s_25s_0_2_6), 
           .COUT(co_mult_29s_25s_0_2_7), .S0(s_mult_29s_25s_0_2_21), .S1(s_mult_29s_25s_0_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_8 (.A0(mult_29s_25s_0_pp_4_23), .A1(mult_29s_25s_0_pp_4_24), 
           .B0(mult_29s_25s_0_pp_5_23), .B1(mult_29s_25s_0_pp_5_24), .CI(co_mult_29s_25s_0_2_7), 
           .COUT(co_mult_29s_25s_0_2_8), .S0(s_mult_29s_25s_0_2_23), .S1(s_mult_29s_25s_0_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_9 (.A0(mult_29s_25s_0_pp_4_25), .A1(mult_29s_25s_0_pp_4_26), 
           .B0(mult_29s_25s_0_pp_5_25), .B1(mult_29s_25s_0_pp_5_26), .CI(co_mult_29s_25s_0_2_8), 
           .COUT(co_mult_29s_25s_0_2_9), .S0(s_mult_29s_25s_0_2_25), .S1(s_mult_29s_25s_0_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_10 (.A0(mult_29s_25s_0_pp_4_27), .A1(mult_29s_25s_0_pp_4_28), 
           .B0(mult_29s_25s_0_pp_5_27), .B1(mult_29s_25s_0_pp_5_28), .CI(co_mult_29s_25s_0_2_9), 
           .S0(s_mult_29s_25s_0_2_27), .S1(s_mult_29s_25s_0_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 mux_237_i6_3_lut_4_lut_3_lut (.A(n30_adj_2140), .B(n1307[15]), 
         .C(n2261[5]), .Z(n1443[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[25:42])
    defparam mux_237_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FADD2B Cadd_mult_29s_25s_0_3_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_6_14), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_7_14), .CI(GND_net), .COUT(co_mult_29s_25s_0_3_1), 
           .S1(s_mult_29s_25s_0_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_2 (.A0(mult_29s_25s_0_pp_6_15), .A1(mult_29s_25s_0_pp_6_16), 
           .B0(mult_29s_25s_0_pp_7_15), .B1(mult_29s_25s_0_pp_7_16), .CI(co_mult_29s_25s_0_3_1), 
           .COUT(co_mult_29s_25s_0_3_2), .S0(s_mult_29s_25s_0_3_15), .S1(s_mult_29s_25s_0_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_3 (.A0(mult_29s_25s_0_pp_6_17), .A1(mult_29s_25s_0_pp_6_18), 
           .B0(mult_29s_25s_0_pp_7_17), .B1(mult_29s_25s_0_pp_7_18), .CI(co_mult_29s_25s_0_3_2), 
           .COUT(co_mult_29s_25s_0_3_3), .S0(s_mult_29s_25s_0_3_17), .S1(s_mult_29s_25s_0_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_4 (.A0(mult_29s_25s_0_pp_6_19), .A1(mult_29s_25s_0_pp_6_20), 
           .B0(mult_29s_25s_0_pp_7_19), .B1(mult_29s_25s_0_pp_7_20), .CI(co_mult_29s_25s_0_3_3), 
           .COUT(co_mult_29s_25s_0_3_4), .S0(s_mult_29s_25s_0_3_19), .S1(s_mult_29s_25s_0_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_5 (.A0(mult_29s_25s_0_pp_6_21), .A1(mult_29s_25s_0_pp_6_22), 
           .B0(mult_29s_25s_0_pp_7_21), .B1(mult_29s_25s_0_pp_7_22), .CI(co_mult_29s_25s_0_3_4), 
           .COUT(co_mult_29s_25s_0_3_5), .S0(s_mult_29s_25s_0_3_21), .S1(s_mult_29s_25s_0_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_6 (.A0(mult_29s_25s_0_pp_6_23), .A1(mult_29s_25s_0_pp_6_24), 
           .B0(mult_29s_25s_0_pp_7_23), .B1(mult_29s_25s_0_pp_7_24), .CI(co_mult_29s_25s_0_3_5), 
           .COUT(co_mult_29s_25s_0_3_6), .S0(s_mult_29s_25s_0_3_23), .S1(s_mult_29s_25s_0_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_7 (.A0(mult_29s_25s_0_pp_6_25), .A1(mult_29s_25s_0_pp_6_26), 
           .B0(mult_29s_25s_0_pp_7_25), .B1(mult_29s_25s_0_pp_7_26), .CI(co_mult_29s_25s_0_3_6), 
           .COUT(co_mult_29s_25s_0_3_7), .S0(s_mult_29s_25s_0_3_25), .S1(s_mult_29s_25s_0_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_8 (.A0(mult_29s_25s_0_pp_6_27), .A1(mult_29s_25s_0_pp_6_28), 
           .B0(mult_29s_25s_0_pp_7_27), .B1(mult_29s_25s_0_pp_7_28), .CI(co_mult_29s_25s_0_3_7), 
           .S0(s_mult_29s_25s_0_3_27), .S1(s_mult_29s_25s_0_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_4_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_8_18), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_9_18), .CI(GND_net), .COUT(co_mult_29s_25s_0_4_1), 
           .S1(s_mult_29s_25s_0_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_2 (.A0(mult_29s_25s_0_pp_8_19), .A1(mult_29s_25s_0_pp_8_20), 
           .B0(mult_29s_25s_0_pp_9_19), .B1(mult_29s_25s_0_pp_9_20), .CI(co_mult_29s_25s_0_4_1), 
           .COUT(co_mult_29s_25s_0_4_2), .S0(s_mult_29s_25s_0_4_19), .S1(s_mult_29s_25s_0_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_3 (.A0(mult_29s_25s_0_pp_8_21), .A1(mult_29s_25s_0_pp_8_22), 
           .B0(mult_29s_25s_0_pp_9_21), .B1(mult_29s_25s_0_pp_9_22), .CI(co_mult_29s_25s_0_4_2), 
           .COUT(co_mult_29s_25s_0_4_3), .S0(s_mult_29s_25s_0_4_21), .S1(s_mult_29s_25s_0_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_4 (.A0(mult_29s_25s_0_pp_8_23), .A1(mult_29s_25s_0_pp_8_24), 
           .B0(mult_29s_25s_0_pp_9_23), .B1(mult_29s_25s_0_pp_9_24), .CI(co_mult_29s_25s_0_4_3), 
           .COUT(co_mult_29s_25s_0_4_4), .S0(s_mult_29s_25s_0_4_23), .S1(s_mult_29s_25s_0_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_5 (.A0(mult_29s_25s_0_pp_8_25), .A1(mult_29s_25s_0_pp_8_26), 
           .B0(mult_29s_25s_0_pp_9_25), .B1(mult_29s_25s_0_pp_9_26), .CI(co_mult_29s_25s_0_4_4), 
           .COUT(co_mult_29s_25s_0_4_5), .S0(s_mult_29s_25s_0_4_25), .S1(s_mult_29s_25s_0_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_6 (.A0(mult_29s_25s_0_pp_8_27), .A1(mult_29s_25s_0_pp_8_28), 
           .B0(mult_29s_25s_0_pp_9_27), .B1(mult_29s_25s_0_pp_9_28), .CI(co_mult_29s_25s_0_4_5), 
           .S0(s_mult_29s_25s_0_4_27), .S1(s_mult_29s_25s_0_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_5_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_10_22), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_11_22), .CI(GND_net), .COUT(co_mult_29s_25s_0_5_1), 
           .S1(s_mult_29s_25s_0_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_2 (.A0(mult_29s_25s_0_pp_10_23), .A1(mult_29s_25s_0_pp_10_24), 
           .B0(mult_29s_25s_0_pp_11_23), .B1(mult_29s_25s_0_pp_11_24), .CI(co_mult_29s_25s_0_5_1), 
           .COUT(co_mult_29s_25s_0_5_2), .S0(s_mult_29s_25s_0_5_23), .S1(s_mult_29s_25s_0_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_3 (.A0(mult_29s_25s_0_pp_10_25), .A1(mult_29s_25s_0_pp_10_26), 
           .B0(mult_29s_25s_0_pp_11_25), .B1(mult_29s_25s_0_pp_11_26), .CI(co_mult_29s_25s_0_5_2), 
           .COUT(co_mult_29s_25s_0_5_3), .S0(s_mult_29s_25s_0_5_25), .S1(s_mult_29s_25s_0_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_4 (.A0(mult_29s_25s_0_pp_10_27), .A1(mult_29s_25s_0_pp_10_28), 
           .B0(mult_29s_25s_0_pp_11_27), .B1(mult_29s_25s_0_pp_11_28), .CI(co_mult_29s_25s_0_5_3), 
           .S0(s_mult_29s_25s_0_5_27), .S1(s_mult_29s_25s_0_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 mux_135_i22_4_lut (.A(backOut2[21]), .B(backOut3[21]), .C(n21321), 
         .D(n9), .Z(n551[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i22_4_lut.init = 16'h0aca;
    FADD2B Cadd_mult_29s_25s_0_6_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_12_24), 
           .B0(GND_net), .B1(VCC_net), .CI(GND_net), .COUT(co_mult_29s_25s_0_6_1), 
           .S1(s_mult_29s_25s_0_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_2 (.A0(mult_29s_25s_0_pp_12_25), .A1(mult_29s_25s_0_pp_12_26), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_1), .COUT(co_mult_29s_25s_0_6_2), 
           .S0(s_mult_29s_25s_0_6_25), .S1(s_mult_29s_25s_0_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_3 (.A0(mult_29s_25s_0_pp_12_27), .A1(mult_29s_25s_0_pp_12_28), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_2), .S0(s_mult_29s_25s_0_6_27), 
           .S1(s_mult_29s_25s_0_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_7_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_0_4), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_2_4), .CI(GND_net), .COUT(co_mult_29s_25s_0_7_1), 
           .S1(multOut_28__N_1217[4])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_2 (.A0(s_mult_29s_25s_0_0_5), .A1(s_mult_29s_25s_0_0_6), 
           .B0(mult_29s_25s_0_pp_2_5), .B1(s_mult_29s_25s_0_1_6), .CI(co_mult_29s_25s_0_7_1), 
           .COUT(co_mult_29s_25s_0_7_2), .S0(multOut_28__N_1217[5]), .S1(multOut_28__N_1217[6])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_3 (.A0(s_mult_29s_25s_0_0_7), .A1(s_mult_29s_25s_0_0_8), 
           .B0(s_mult_29s_25s_0_1_7), .B1(s_mult_29s_25s_0_1_8), .CI(co_mult_29s_25s_0_7_2), 
           .COUT(co_mult_29s_25s_0_7_3), .S0(multOut_28__N_1217[7]), .S1(s_mult_29s_25s_0_7_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_4 (.A0(s_mult_29s_25s_0_0_9), .A1(s_mult_29s_25s_0_0_10), 
           .B0(s_mult_29s_25s_0_1_9), .B1(s_mult_29s_25s_0_1_10), .CI(co_mult_29s_25s_0_7_3), 
           .COUT(co_mult_29s_25s_0_7_4), .S0(s_mult_29s_25s_0_7_9), .S1(s_mult_29s_25s_0_7_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_5 (.A0(s_mult_29s_25s_0_0_11), .A1(s_mult_29s_25s_0_0_12), 
           .B0(s_mult_29s_25s_0_1_11), .B1(s_mult_29s_25s_0_1_12), .CI(co_mult_29s_25s_0_7_4), 
           .COUT(co_mult_29s_25s_0_7_5), .S0(s_mult_29s_25s_0_7_11), .S1(s_mult_29s_25s_0_7_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_6 (.A0(s_mult_29s_25s_0_0_13), .A1(s_mult_29s_25s_0_0_14), 
           .B0(s_mult_29s_25s_0_1_13), .B1(s_mult_29s_25s_0_1_14), .CI(co_mult_29s_25s_0_7_5), 
           .COUT(co_mult_29s_25s_0_7_6), .S0(s_mult_29s_25s_0_7_13), .S1(s_mult_29s_25s_0_7_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_7 (.A0(s_mult_29s_25s_0_0_15), .A1(s_mult_29s_25s_0_0_16), 
           .B0(s_mult_29s_25s_0_1_15), .B1(s_mult_29s_25s_0_1_16), .CI(co_mult_29s_25s_0_7_6), 
           .COUT(co_mult_29s_25s_0_7_7), .S0(s_mult_29s_25s_0_7_15), .S1(s_mult_29s_25s_0_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_8 (.A0(s_mult_29s_25s_0_0_17), .A1(s_mult_29s_25s_0_0_18), 
           .B0(s_mult_29s_25s_0_1_17), .B1(s_mult_29s_25s_0_1_18), .CI(co_mult_29s_25s_0_7_7), 
           .COUT(co_mult_29s_25s_0_7_8), .S0(s_mult_29s_25s_0_7_17), .S1(s_mult_29s_25s_0_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_9 (.A0(s_mult_29s_25s_0_0_19), .A1(s_mult_29s_25s_0_0_20), 
           .B0(s_mult_29s_25s_0_1_19), .B1(s_mult_29s_25s_0_1_20), .CI(co_mult_29s_25s_0_7_8), 
           .COUT(co_mult_29s_25s_0_7_9), .S0(s_mult_29s_25s_0_7_19), .S1(s_mult_29s_25s_0_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_10 (.A0(s_mult_29s_25s_0_0_21), .A1(s_mult_29s_25s_0_0_22), 
           .B0(s_mult_29s_25s_0_1_21), .B1(s_mult_29s_25s_0_1_22), .CI(co_mult_29s_25s_0_7_9), 
           .COUT(co_mult_29s_25s_0_7_10), .S0(s_mult_29s_25s_0_7_21), .S1(s_mult_29s_25s_0_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_11 (.A0(s_mult_29s_25s_0_0_23), .A1(s_mult_29s_25s_0_0_24), 
           .B0(s_mult_29s_25s_0_1_23), .B1(s_mult_29s_25s_0_1_24), .CI(co_mult_29s_25s_0_7_10), 
           .COUT(co_mult_29s_25s_0_7_11), .S0(s_mult_29s_25s_0_7_23), .S1(s_mult_29s_25s_0_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_12 (.A0(s_mult_29s_25s_0_0_25), .A1(s_mult_29s_25s_0_0_26), 
           .B0(s_mult_29s_25s_0_1_25), .B1(s_mult_29s_25s_0_1_26), .CI(co_mult_29s_25s_0_7_11), 
           .COUT(co_mult_29s_25s_0_7_12), .S0(s_mult_29s_25s_0_7_25), .S1(s_mult_29s_25s_0_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_13 (.A0(s_mult_29s_25s_0_0_27), .A1(s_mult_29s_25s_0_0_28), 
           .B0(s_mult_29s_25s_0_1_27), .B1(s_mult_29s_25s_0_1_28), .CI(co_mult_29s_25s_0_7_12), 
           .S0(s_mult_29s_25s_0_7_27), .S1(s_mult_29s_25s_0_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_8_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_2_12), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_6_12), .CI(GND_net), .COUT(co_mult_29s_25s_0_8_1), 
           .S1(s_mult_29s_25s_0_8_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_2 (.A0(s_mult_29s_25s_0_2_13), .A1(s_mult_29s_25s_0_2_14), 
           .B0(mult_29s_25s_0_pp_6_13), .B1(s_mult_29s_25s_0_3_14), .CI(co_mult_29s_25s_0_8_1), 
           .COUT(co_mult_29s_25s_0_8_2), .S0(s_mult_29s_25s_0_8_13), .S1(s_mult_29s_25s_0_8_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_3 (.A0(s_mult_29s_25s_0_2_15), .A1(s_mult_29s_25s_0_2_16), 
           .B0(s_mult_29s_25s_0_3_15), .B1(s_mult_29s_25s_0_3_16), .CI(co_mult_29s_25s_0_8_2), 
           .COUT(co_mult_29s_25s_0_8_3), .S0(s_mult_29s_25s_0_8_15), .S1(s_mult_29s_25s_0_8_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_4 (.A0(s_mult_29s_25s_0_2_17), .A1(s_mult_29s_25s_0_2_18), 
           .B0(s_mult_29s_25s_0_3_17), .B1(s_mult_29s_25s_0_3_18), .CI(co_mult_29s_25s_0_8_3), 
           .COUT(co_mult_29s_25s_0_8_4), .S0(s_mult_29s_25s_0_8_17), .S1(s_mult_29s_25s_0_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_5 (.A0(s_mult_29s_25s_0_2_19), .A1(s_mult_29s_25s_0_2_20), 
           .B0(s_mult_29s_25s_0_3_19), .B1(s_mult_29s_25s_0_3_20), .CI(co_mult_29s_25s_0_8_4), 
           .COUT(co_mult_29s_25s_0_8_5), .S0(s_mult_29s_25s_0_8_19), .S1(s_mult_29s_25s_0_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_6 (.A0(s_mult_29s_25s_0_2_21), .A1(s_mult_29s_25s_0_2_22), 
           .B0(s_mult_29s_25s_0_3_21), .B1(s_mult_29s_25s_0_3_22), .CI(co_mult_29s_25s_0_8_5), 
           .COUT(co_mult_29s_25s_0_8_6), .S0(s_mult_29s_25s_0_8_21), .S1(s_mult_29s_25s_0_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_7 (.A0(s_mult_29s_25s_0_2_23), .A1(s_mult_29s_25s_0_2_24), 
           .B0(s_mult_29s_25s_0_3_23), .B1(s_mult_29s_25s_0_3_24), .CI(co_mult_29s_25s_0_8_6), 
           .COUT(co_mult_29s_25s_0_8_7), .S0(s_mult_29s_25s_0_8_23), .S1(s_mult_29s_25s_0_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_8 (.A0(s_mult_29s_25s_0_2_25), .A1(s_mult_29s_25s_0_2_26), 
           .B0(s_mult_29s_25s_0_3_25), .B1(s_mult_29s_25s_0_3_26), .CI(co_mult_29s_25s_0_8_7), 
           .COUT(co_mult_29s_25s_0_8_8), .S0(s_mult_29s_25s_0_8_25), .S1(s_mult_29s_25s_0_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_9 (.A0(s_mult_29s_25s_0_2_27), .A1(s_mult_29s_25s_0_2_28), 
           .B0(s_mult_29s_25s_0_3_27), .B1(s_mult_29s_25s_0_3_28), .CI(co_mult_29s_25s_0_8_8), 
           .S0(s_mult_29s_25s_0_8_27), .S1(s_mult_29s_25s_0_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_9_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_4_20), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_10_20), .CI(GND_net), .COUT(co_mult_29s_25s_0_9_1), 
           .S1(s_mult_29s_25s_0_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_2 (.A0(s_mult_29s_25s_0_4_21), .A1(s_mult_29s_25s_0_4_22), 
           .B0(mult_29s_25s_0_pp_10_21), .B1(s_mult_29s_25s_0_5_22), .CI(co_mult_29s_25s_0_9_1), 
           .COUT(co_mult_29s_25s_0_9_2), .S0(s_mult_29s_25s_0_9_21), .S1(s_mult_29s_25s_0_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_3 (.A0(s_mult_29s_25s_0_4_23), .A1(s_mult_29s_25s_0_4_24), 
           .B0(s_mult_29s_25s_0_5_23), .B1(s_mult_29s_25s_0_5_24), .CI(co_mult_29s_25s_0_9_2), 
           .COUT(co_mult_29s_25s_0_9_3), .S0(s_mult_29s_25s_0_9_23), .S1(s_mult_29s_25s_0_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_4 (.A0(s_mult_29s_25s_0_4_25), .A1(s_mult_29s_25s_0_4_26), 
           .B0(s_mult_29s_25s_0_5_25), .B1(s_mult_29s_25s_0_5_26), .CI(co_mult_29s_25s_0_9_3), 
           .COUT(co_mult_29s_25s_0_9_4), .S0(s_mult_29s_25s_0_9_25), .S1(s_mult_29s_25s_0_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_5 (.A0(s_mult_29s_25s_0_4_27), .A1(s_mult_29s_25s_0_4_28), 
           .B0(s_mult_29s_25s_0_5_27), .B1(s_mult_29s_25s_0_5_28), .CI(co_mult_29s_25s_0_9_4), 
           .S0(s_mult_29s_25s_0_9_27), .S1(s_mult_29s_25s_0_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 mux_244_i9_3_lut_4_lut_3_lut (.A(n30_adj_2141), .B(n1328[15]), 
         .C(n2273[8]), .Z(n1487[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(362[25:42])
    defparam mux_244_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FADD2B Cadd_mult_29s_25s_0_10_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_7_8), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_4_8), .CI(GND_net), .COUT(co_mult_29s_25s_0_10_1), 
           .S1(multOut_28__N_1217[8])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_2 (.A0(s_mult_29s_25s_0_7_9), .A1(s_mult_29s_25s_0_7_10), 
           .B0(mult_29s_25s_0_pp_4_9), .B1(s_mult_29s_25s_0_2_10), .CI(co_mult_29s_25s_0_10_1), 
           .COUT(co_mult_29s_25s_0_10_2), .S0(multOut_28__N_1217[9]), .S1(multOut_28__N_1217[10])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_3 (.A0(s_mult_29s_25s_0_7_11), .A1(s_mult_29s_25s_0_7_12), 
           .B0(s_mult_29s_25s_0_2_11), .B1(s_mult_29s_25s_0_8_12), .CI(co_mult_29s_25s_0_10_2), 
           .COUT(co_mult_29s_25s_0_10_3), .S0(multOut_28__N_1217[11]), .S1(multOut_28__N_1217[12])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_4 (.A0(s_mult_29s_25s_0_7_13), .A1(s_mult_29s_25s_0_7_14), 
           .B0(s_mult_29s_25s_0_8_13), .B1(s_mult_29s_25s_0_8_14), .CI(co_mult_29s_25s_0_10_3), 
           .COUT(co_mult_29s_25s_0_10_4), .S0(multOut_28__N_1217[13]), .S1(multOut_28__N_1217[14])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_5 (.A0(s_mult_29s_25s_0_7_15), .A1(s_mult_29s_25s_0_7_16), 
           .B0(s_mult_29s_25s_0_8_15), .B1(s_mult_29s_25s_0_8_16), .CI(co_mult_29s_25s_0_10_4), 
           .COUT(co_mult_29s_25s_0_10_5), .S0(multOut_28__N_1217[15]), .S1(s_mult_29s_25s_0_10_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_6 (.A0(s_mult_29s_25s_0_7_17), .A1(s_mult_29s_25s_0_7_18), 
           .B0(s_mult_29s_25s_0_8_17), .B1(s_mult_29s_25s_0_8_18), .CI(co_mult_29s_25s_0_10_5), 
           .COUT(co_mult_29s_25s_0_10_6), .S0(s_mult_29s_25s_0_10_17), .S1(s_mult_29s_25s_0_10_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_7 (.A0(s_mult_29s_25s_0_7_19), .A1(s_mult_29s_25s_0_7_20), 
           .B0(s_mult_29s_25s_0_8_19), .B1(s_mult_29s_25s_0_8_20), .CI(co_mult_29s_25s_0_10_6), 
           .COUT(co_mult_29s_25s_0_10_7), .S0(s_mult_29s_25s_0_10_19), .S1(s_mult_29s_25s_0_10_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_8 (.A0(s_mult_29s_25s_0_7_21), .A1(s_mult_29s_25s_0_7_22), 
           .B0(s_mult_29s_25s_0_8_21), .B1(s_mult_29s_25s_0_8_22), .CI(co_mult_29s_25s_0_10_7), 
           .COUT(co_mult_29s_25s_0_10_8), .S0(s_mult_29s_25s_0_10_21), .S1(s_mult_29s_25s_0_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_9 (.A0(s_mult_29s_25s_0_7_23), .A1(s_mult_29s_25s_0_7_24), 
           .B0(s_mult_29s_25s_0_8_23), .B1(s_mult_29s_25s_0_8_24), .CI(co_mult_29s_25s_0_10_8), 
           .COUT(co_mult_29s_25s_0_10_9), .S0(s_mult_29s_25s_0_10_23), .S1(s_mult_29s_25s_0_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_10 (.A0(s_mult_29s_25s_0_7_25), .A1(s_mult_29s_25s_0_7_26), 
           .B0(s_mult_29s_25s_0_8_25), .B1(s_mult_29s_25s_0_8_26), .CI(co_mult_29s_25s_0_10_9), 
           .COUT(co_mult_29s_25s_0_10_10), .S0(s_mult_29s_25s_0_10_25), 
           .S1(s_mult_29s_25s_0_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_11 (.A0(s_mult_29s_25s_0_7_27), .A1(s_mult_29s_25s_0_7_28), 
           .B0(s_mult_29s_25s_0_8_27), .B1(s_mult_29s_25s_0_8_28), .CI(co_mult_29s_25s_0_10_10), 
           .S0(s_mult_29s_25s_0_10_27), .S1(s_mult_29s_25s_0_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_11_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_9_24), 
           .B0(GND_net), .B1(s_mult_29s_25s_0_6_24), .CI(GND_net), .COUT(co_mult_29s_25s_0_11_1), 
           .S1(s_mult_29s_25s_0_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_2 (.A0(s_mult_29s_25s_0_9_25), .A1(s_mult_29s_25s_0_9_26), 
           .B0(s_mult_29s_25s_0_6_25), .B1(s_mult_29s_25s_0_6_26), .CI(co_mult_29s_25s_0_11_1), 
           .COUT(co_mult_29s_25s_0_11_2), .S0(s_mult_29s_25s_0_11_25), .S1(s_mult_29s_25s_0_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_3 (.A0(s_mult_29s_25s_0_9_27), .A1(s_mult_29s_25s_0_9_28), 
           .B0(s_mult_29s_25s_0_6_27), .B1(s_mult_29s_25s_0_6_28), .CI(co_mult_29s_25s_0_11_2), 
           .S0(s_mult_29s_25s_0_11_27), .S1(s_mult_29s_25s_0_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 mux_244_i10_3_lut_4_lut_3_lut (.A(n30_adj_2141), .B(n1328[15]), 
         .C(n2273[9]), .Z(n1487[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(362[25:42])
    defparam mux_244_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FADD2B Cadd_t_mult_29s_25s_0_12_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_10_16), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_8_16), .CI(GND_net), .COUT(co_t_mult_29s_25s_0_12_1), 
           .S1(multOut_28__N_1217[16])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_2 (.A0(s_mult_29s_25s_0_10_17), .A1(s_mult_29s_25s_0_10_18), 
           .B0(mult_29s_25s_0_pp_8_17), .B1(s_mult_29s_25s_0_4_18), .CI(co_t_mult_29s_25s_0_12_1), 
           .COUT(co_t_mult_29s_25s_0_12_2), .S0(multOut_28__N_1217[17]), 
           .S1(multOut_28__N_1217[18])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_3 (.A0(s_mult_29s_25s_0_10_19), .A1(s_mult_29s_25s_0_10_20), 
           .B0(s_mult_29s_25s_0_4_19), .B1(s_mult_29s_25s_0_9_20), .CI(co_t_mult_29s_25s_0_12_2), 
           .COUT(co_t_mult_29s_25s_0_12_3), .S0(multOut_28__N_1217[19]), 
           .S1(multOut_28__N_1217[20])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_4 (.A0(s_mult_29s_25s_0_10_21), .A1(s_mult_29s_25s_0_10_22), 
           .B0(s_mult_29s_25s_0_9_21), .B1(s_mult_29s_25s_0_9_22), .CI(co_t_mult_29s_25s_0_12_3), 
           .COUT(co_t_mult_29s_25s_0_12_4), .S0(multOut_28__N_1217[21]), 
           .S1(multOut_28__N_1217[22])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_5 (.A0(s_mult_29s_25s_0_10_23), .A1(s_mult_29s_25s_0_10_24), 
           .B0(s_mult_29s_25s_0_9_23), .B1(s_mult_29s_25s_0_11_24), .CI(co_t_mult_29s_25s_0_12_4), 
           .COUT(co_t_mult_29s_25s_0_12_5), .S0(multOut_28__N_1217[23]), 
           .S1(multOut_28__N_1217[24])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_6 (.A0(s_mult_29s_25s_0_10_25), .A1(s_mult_29s_25s_0_10_26), 
           .B0(s_mult_29s_25s_0_11_25), .B1(s_mult_29s_25s_0_11_26), .CI(co_t_mult_29s_25s_0_12_5), 
           .COUT(co_t_mult_29s_25s_0_12_6), .S0(multOut_28__N_1217[25]), 
           .S1(multOut_28__N_1217[26])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_7 (.A0(s_mult_29s_25s_0_10_27), .A1(s_mult_29s_25s_0_10_28), 
           .B0(s_mult_29s_25s_0_11_27), .B1(s_mult_29s_25s_0_11_28), .CI(co_t_mult_29s_25s_0_12_6), 
           .S0(multOut_28__N_1217[27]), .S1(multOut_28__N_1217[28])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_0), .CO(mco), .P0(multOut_28__N_1217[1]), 
          .P1(mult_29s_25s_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco), .CO(mco_1), .P0(mult_29s_25s_0_pp_0_3), 
          .P1(mult_29s_25s_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_1), .CO(mco_2), .P0(mult_29s_25s_0_pp_0_5), 
          .P1(mult_29s_25s_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_2), .CO(mco_3), .P0(mult_29s_25s_0_pp_0_7), 
          .P1(mult_29s_25s_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_3), .CO(mco_4), .P0(mult_29s_25s_0_pp_0_9), 
          .P1(mult_29s_25s_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_4), .CO(mco_5), .P0(mult_29s_25s_0_pp_0_11), 
          .P1(mult_29s_25s_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_5), .CO(mco_6), .P0(mult_29s_25s_0_pp_0_13), 
          .P1(mult_29s_25s_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_6), .CO(mco_7), .P0(mult_29s_25s_0_pp_0_15), 
          .P1(mult_29s_25s_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_7), .CO(mco_8), .P0(mult_29s_25s_0_pp_0_17), 
          .P1(mult_29s_25s_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_8), .CO(mco_9), .P0(mult_29s_25s_0_pp_0_19), 
          .P1(mult_29s_25s_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_9), .CO(mco_10), .P0(mult_29s_25s_0_pp_0_21), 
          .P1(mult_29s_25s_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_10), .CO(mco_11), .P0(mult_29s_25s_0_pp_0_23), 
          .P1(mult_29s_25s_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_11), .CO(mco_12), .P0(mult_29s_25s_0_pp_0_25), 
          .P1(mult_29s_25s_0_pp_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_13 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_12), .P0(mult_29s_25s_0_pp_0_27), .P1(mult_29s_25s_0_pp_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_2), .CO(mco_14), 
          .P0(mult_29s_25s_0_pp_1_3), .P1(mult_29s_25s_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_14), .CO(mco_15), .P0(mult_29s_25s_0_pp_1_5), 
          .P1(mult_29s_25s_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_15), .CO(mco_16), .P0(mult_29s_25s_0_pp_1_7), 
          .P1(mult_29s_25s_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_16), .CO(mco_17), .P0(mult_29s_25s_0_pp_1_9), 
          .P1(mult_29s_25s_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_17), .CO(mco_18), .P0(mult_29s_25s_0_pp_1_11), 
          .P1(mult_29s_25s_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_18), .CO(mco_19), .P0(mult_29s_25s_0_pp_1_13), 
          .P1(mult_29s_25s_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_19), .CO(mco_20), .P0(mult_29s_25s_0_pp_1_15), 
          .P1(mult_29s_25s_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_20), .CO(mco_21), .P0(mult_29s_25s_0_pp_1_17), 
          .P1(mult_29s_25s_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_21), .CO(mco_22), .P0(mult_29s_25s_0_pp_1_19), 
          .P1(mult_29s_25s_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_22), .CO(mco_23), .P0(mult_29s_25s_0_pp_1_21), 
          .P1(mult_29s_25s_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_23), .CO(mco_24), .P0(mult_29s_25s_0_pp_1_23), 
          .P1(mult_29s_25s_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_24), .CO(mco_25), .P0(mult_29s_25s_0_pp_1_25), 
          .P1(mult_29s_25s_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_25), .P0(mult_29s_25s_0_pp_1_27), .P1(mult_29s_25s_0_pp_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_4), .CO(mco_28), 
          .P0(mult_29s_25s_0_pp_2_5), .P1(mult_29s_25s_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_28), .CO(mco_29), .P0(mult_29s_25s_0_pp_2_7), 
          .P1(mult_29s_25s_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_29), .CO(mco_30), .P0(mult_29s_25s_0_pp_2_9), 
          .P1(mult_29s_25s_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_30), .CO(mco_31), .P0(mult_29s_25s_0_pp_2_11), 
          .P1(mult_29s_25s_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_31), .CO(mco_32), .P0(mult_29s_25s_0_pp_2_13), 
          .P1(mult_29s_25s_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_32), .CO(mco_33), .P0(mult_29s_25s_0_pp_2_15), 
          .P1(mult_29s_25s_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_33), .CO(mco_34), .P0(mult_29s_25s_0_pp_2_17), 
          .P1(mult_29s_25s_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_34), .CO(mco_35), .P0(mult_29s_25s_0_pp_2_19), 
          .P1(mult_29s_25s_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_35), .CO(mco_36), .P0(mult_29s_25s_0_pp_2_21), 
          .P1(mult_29s_25s_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_36), .CO(mco_37), .P0(mult_29s_25s_0_pp_2_23), 
          .P1(mult_29s_25s_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_37), .CO(mco_38), .P0(mult_29s_25s_0_pp_2_25), 
          .P1(mult_29s_25s_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_38), .P0(mult_29s_25s_0_pp_2_27), .P1(mult_29s_25s_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_6), .CO(mco_42), 
          .P0(mult_29s_25s_0_pp_3_7), .P1(mult_29s_25s_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_42), .CO(mco_43), .P0(mult_29s_25s_0_pp_3_9), 
          .P1(mult_29s_25s_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_43), .CO(mco_44), .P0(mult_29s_25s_0_pp_3_11), 
          .P1(mult_29s_25s_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_44), .CO(mco_45), .P0(mult_29s_25s_0_pp_3_13), 
          .P1(mult_29s_25s_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_45), .CO(mco_46), .P0(mult_29s_25s_0_pp_3_15), 
          .P1(mult_29s_25s_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_46), .CO(mco_47), .P0(mult_29s_25s_0_pp_3_17), 
          .P1(mult_29s_25s_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_47), .CO(mco_48), .P0(mult_29s_25s_0_pp_3_19), 
          .P1(mult_29s_25s_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_48), .CO(mco_49), .P0(mult_29s_25s_0_pp_3_21), 
          .P1(mult_29s_25s_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_49), .CO(mco_50), .P0(mult_29s_25s_0_pp_3_23), 
          .P1(mult_29s_25s_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_50), .CO(mco_51), .P0(mult_29s_25s_0_pp_3_25), 
          .P1(mult_29s_25s_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[4]), .B1(multIn2[4]), .B2(multIn2[4]), 
          .B3(multIn2[4]), .CI(mco_51), .P0(mult_29s_25s_0_pp_3_27), .P1(mult_29s_25s_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mult_29s_25s_0_cin_lr_8), .CO(mco_56), 
          .P0(mult_29s_25s_0_pp_4_9), .P1(mult_29s_25s_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_56), .CO(mco_57), .P0(mult_29s_25s_0_pp_4_11), 
          .P1(mult_29s_25s_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_57), .CO(mco_58), .P0(mult_29s_25s_0_pp_4_13), 
          .P1(mult_29s_25s_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_58), .CO(mco_59), .P0(mult_29s_25s_0_pp_4_15), 
          .P1(mult_29s_25s_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_59), .CO(mco_60), .P0(mult_29s_25s_0_pp_4_17), 
          .P1(mult_29s_25s_0_pp_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_60), .CO(mco_61), .P0(mult_29s_25s_0_pp_4_19), 
          .P1(mult_29s_25s_0_pp_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_61), .CO(mco_62), .P0(mult_29s_25s_0_pp_4_21), 
          .P1(mult_29s_25s_0_pp_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_62), .CO(mco_63), .P0(mult_29s_25s_0_pp_4_23), 
          .P1(mult_29s_25s_0_pp_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_63), .CO(mco_64), .P0(mult_29s_25s_0_pp_4_25), 
          .P1(mult_29s_25s_0_pp_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(multIn2[4]), .B2(GND_net), 
          .B3(multIn2[4]), .CI(mco_64), .P0(mult_29s_25s_0_pp_4_27), .P1(mult_29s_25s_0_pp_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_10), .CO(mco_70), .P0(mult_29s_25s_0_pp_5_11), 
          .P1(mult_29s_25s_0_pp_5_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_70), .CO(mco_71), .P0(mult_29s_25s_0_pp_5_13), 
          .P1(mult_29s_25s_0_pp_5_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_71), .CO(mco_72), .P0(mult_29s_25s_0_pp_5_15), 
          .P1(mult_29s_25s_0_pp_5_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_72), .CO(mco_73), .P0(mult_29s_25s_0_pp_5_17), 
          .P1(mult_29s_25s_0_pp_5_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_73), .CO(mco_74), .P0(mult_29s_25s_0_pp_5_19), 
          .P1(mult_29s_25s_0_pp_5_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_74), .CO(mco_75), .P0(mult_29s_25s_0_pp_5_21), 
          .P1(mult_29s_25s_0_pp_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_75), .CO(mco_76), .P0(mult_29s_25s_0_pp_5_23), 
          .P1(mult_29s_25s_0_pp_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_76), .CO(mco_77), .P0(mult_29s_25s_0_pp_5_25), 
          .P1(mult_29s_25s_0_pp_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_77), .P0(mult_29s_25s_0_pp_5_27), .P1(mult_29s_25s_0_pp_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_12), .CO(mco_84), .P0(mult_29s_25s_0_pp_6_13), 
          .P1(mult_29s_25s_0_pp_6_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_84), .CO(mco_85), .P0(mult_29s_25s_0_pp_6_15), 
          .P1(mult_29s_25s_0_pp_6_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_85), .CO(mco_86), .P0(mult_29s_25s_0_pp_6_17), 
          .P1(mult_29s_25s_0_pp_6_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_86), .CO(mco_87), .P0(mult_29s_25s_0_pp_6_19), 
          .P1(mult_29s_25s_0_pp_6_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_87), .CO(mco_88), .P0(mult_29s_25s_0_pp_6_21), 
          .P1(mult_29s_25s_0_pp_6_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_88), .CO(mco_89), .P0(mult_29s_25s_0_pp_6_23), 
          .P1(mult_29s_25s_0_pp_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_89), .CO(mco_90), .P0(mult_29s_25s_0_pp_6_25), 
          .P1(mult_29s_25s_0_pp_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_90), .P0(mult_29s_25s_0_pp_6_27), .P1(mult_29s_25s_0_pp_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_14), .CO(mco_98), .P0(mult_29s_25s_0_pp_7_15), 
          .P1(mult_29s_25s_0_pp_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_98), .CO(mco_99), .P0(mult_29s_25s_0_pp_7_17), 
          .P1(mult_29s_25s_0_pp_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_99), .CO(mco_100), .P0(mult_29s_25s_0_pp_7_19), 
          .P1(mult_29s_25s_0_pp_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_100), .CO(mco_101), .P0(mult_29s_25s_0_pp_7_21), 
          .P1(mult_29s_25s_0_pp_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_101), .CO(mco_102), .P0(mult_29s_25s_0_pp_7_23), 
          .P1(mult_29s_25s_0_pp_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_102), .CO(mco_103), .P0(mult_29s_25s_0_pp_7_25), 
          .P1(mult_29s_25s_0_pp_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_103), .P0(mult_29s_25s_0_pp_7_27), .P1(mult_29s_25s_0_pp_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_16), .CO(mco_112), .P0(mult_29s_25s_0_pp_8_17), 
          .P1(mult_29s_25s_0_pp_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_112), .CO(mco_113), .P0(mult_29s_25s_0_pp_8_19), 
          .P1(mult_29s_25s_0_pp_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_113), .CO(mco_114), .P0(mult_29s_25s_0_pp_8_21), 
          .P1(mult_29s_25s_0_pp_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_114), .CO(mco_115), .P0(mult_29s_25s_0_pp_8_23), 
          .P1(mult_29s_25s_0_pp_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_115), .CO(mco_116), .P0(mult_29s_25s_0_pp_8_25), 
          .P1(mult_29s_25s_0_pp_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_116), .P0(mult_29s_25s_0_pp_8_27), .P1(mult_29s_25s_0_pp_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 mux_237_i10_3_lut_4_lut_3_lut (.A(n30_adj_2140), .B(n1307[15]), 
         .C(n2261[9]), .Z(n1443[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[25:42])
    defparam mux_237_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    MULT2 mult_29s_25s_0_mult_18_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_18), .CO(mco_126), .P0(mult_29s_25s_0_pp_9_19), 
          .P1(mult_29s_25s_0_pp_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_126), .CO(mco_127), .P0(mult_29s_25s_0_pp_9_21), 
          .P1(mult_29s_25s_0_pp_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_127), .CO(mco_128), .P0(mult_29s_25s_0_pp_9_23), 
          .P1(mult_29s_25s_0_pp_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_128), .CO(mco_129), .P0(mult_29s_25s_0_pp_9_25), 
          .P1(mult_29s_25s_0_pp_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_129), .P0(mult_29s_25s_0_pp_9_27), .P1(mult_29s_25s_0_pp_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_20), .CO(mco_140), .P0(mult_29s_25s_0_pp_10_21), 
          .P1(mult_29s_25s_0_pp_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_140), .CO(mco_141), .P0(mult_29s_25s_0_pp_10_23), 
          .P1(mult_29s_25s_0_pp_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_141), .CO(mco_142), .P0(mult_29s_25s_0_pp_10_25), 
          .P1(mult_29s_25s_0_pp_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_142), .P0(mult_29s_25s_0_pp_10_27), .P1(mult_29s_25s_0_pp_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_22), .CO(mco_154), .P0(mult_29s_25s_0_pp_11_23), 
          .P1(mult_29s_25s_0_pp_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_154), .CO(mco_155), .P0(mult_29s_25s_0_pp_11_25), 
          .P1(mult_29s_25s_0_pp_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_155), .P0(mult_29s_25s_0_pp_11_27), .P1(mult_29s_25s_0_pp_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    PFUMX i17488 (.BLUT(n22093), .ALUT(n22094), .C0(ss[1]), .Z(n15696));
    LUT4 mux_237_i7_3_lut_4_lut_3_lut (.A(n30_adj_2140), .B(n1307[15]), 
         .C(n2261[6]), .Z(n1443[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[25:42])
    defparam mux_237_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_244_i6_3_lut_4_lut_3_lut (.A(n30_adj_2141), .B(n1328[15]), 
         .C(n2273[5]), .Z(n1487[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(362[25:42])
    defparam mux_244_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i1_4_lut_adj_53 (.A(n3600), .B(n35_adj_2142), .C(n40), .D(n36), 
         .Z(n4_adj_2134)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_53.init = 16'haaa8;
    FD1P3AX backOut0_i0_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_70), 
            .CK(clk_N_683), .Q(backOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i1.GSR = "DISABLED";
    FD1S3AX multOut_i1 (.D(multOut_28__N_1217[1]), .CK(clk_N_683), .Q(multOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i1.GSR = "ENABLED";
    LUT4 mux_244_i4_3_lut_4_lut_3_lut (.A(n30_adj_2141), .B(n1328[15]), 
         .C(n2273[3]), .Z(n1487[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(362[25:42])
    defparam mux_244_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_135_i1_4_lut (.A(backOut2[0]), .B(backOut3[0]), .C(n21321), 
         .D(n9), .Z(n551[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i1_4_lut.init = 16'h0aca;
    LUT4 mux_135_i23_4_lut (.A(backOut2[22]), .B(backOut3[22]), .C(n21321), 
         .D(n9), .Z(n551[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i23_4_lut.init = 16'h0aca;
    LUT4 mux_135_i24_4_lut (.A(backOut2[23]), .B(backOut3[23]), .C(n21321), 
         .D(n9), .Z(n551[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i24_4_lut.init = 16'h0aca;
    LUT4 i2_4_lut_4_lut_rep_404 (.A(n9_adj_2138), .B(n21342), .C(ss[1]), 
         .Z(n22082)) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i2_4_lut_4_lut_rep_404.init = 16'h8a8a;
    FD1S3AX multOut_i2 (.D(multOut_28__N_1217[2]), .CK(clk_N_683), .Q(multOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i2.GSR = "ENABLED";
    FD1S3AX multOut_i3 (.D(multOut_28__N_1217[3]), .CK(clk_N_683), .Q(multOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i3.GSR = "ENABLED";
    FD1S3AX multOut_i4 (.D(multOut_28__N_1217[4]), .CK(clk_N_683), .Q(multOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i4.GSR = "ENABLED";
    FD1S3AX multOut_i5 (.D(multOut_28__N_1217[5]), .CK(clk_N_683), .Q(multOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i5.GSR = "ENABLED";
    FD1S3AX multOut_i6 (.D(multOut_28__N_1217[6]), .CK(clk_N_683), .Q(multOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i6.GSR = "ENABLED";
    FD1S3AX multOut_i7 (.D(multOut_28__N_1217[7]), .CK(clk_N_683), .Q(multOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i7.GSR = "ENABLED";
    FD1S3AX multOut_i8 (.D(multOut_28__N_1217[8]), .CK(clk_N_683), .Q(multOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i8.GSR = "ENABLED";
    FD1S3AX multOut_i9 (.D(multOut_28__N_1217[9]), .CK(clk_N_683), .Q(multOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i9.GSR = "ENABLED";
    FD1S3AX multOut_i10 (.D(multOut_28__N_1217[10]), .CK(clk_N_683), .Q(multOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i10.GSR = "ENABLED";
    FD1S3AX multOut_i11 (.D(multOut_28__N_1217[11]), .CK(clk_N_683), .Q(multOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i11.GSR = "ENABLED";
    FD1S3AX multOut_i12 (.D(multOut_28__N_1217[12]), .CK(clk_N_683), .Q(multOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i12.GSR = "ENABLED";
    FD1S3AX multOut_i13 (.D(multOut_28__N_1217[13]), .CK(clk_N_683), .Q(multOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i13.GSR = "ENABLED";
    FD1S3AX multOut_i14 (.D(multOut_28__N_1217[14]), .CK(clk_N_683), .Q(multOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i14.GSR = "ENABLED";
    FD1S3AX multOut_i15 (.D(multOut_28__N_1217[15]), .CK(clk_N_683), .Q(multOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i15.GSR = "ENABLED";
    FD1S3AX multOut_i16 (.D(multOut_28__N_1217[16]), .CK(clk_N_683), .Q(multOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i16.GSR = "ENABLED";
    FD1S3AX multOut_i17 (.D(multOut_28__N_1217[17]), .CK(clk_N_683), .Q(multOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i17.GSR = "ENABLED";
    FD1S3AX multOut_i18 (.D(multOut_28__N_1217[18]), .CK(clk_N_683), .Q(multOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i18.GSR = "ENABLED";
    FD1S3AX multOut_i19 (.D(multOut_28__N_1217[19]), .CK(clk_N_683), .Q(multOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i19.GSR = "ENABLED";
    FD1S3AX multOut_i20 (.D(multOut_28__N_1217[20]), .CK(clk_N_683), .Q(multOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i20.GSR = "ENABLED";
    FD1S3AX multOut_i21 (.D(multOut_28__N_1217[21]), .CK(clk_N_683), .Q(multOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i21.GSR = "ENABLED";
    FD1S3AX multOut_i22 (.D(multOut_28__N_1217[22]), .CK(clk_N_683), .Q(multOut[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i22.GSR = "ENABLED";
    FD1S3AX multOut_i23 (.D(multOut_28__N_1217[23]), .CK(clk_N_683), .Q(multOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i23.GSR = "ENABLED";
    FD1S3AX multOut_i24 (.D(multOut_28__N_1217[24]), .CK(clk_N_683), .Q(multOut[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i24.GSR = "ENABLED";
    FD1S3AX multOut_i25 (.D(multOut_28__N_1217[25]), .CK(clk_N_683), .Q(multOut[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i25.GSR = "ENABLED";
    FD1S3AX multOut_i26 (.D(multOut_28__N_1217[26]), .CK(clk_N_683), .Q(multOut[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i26.GSR = "ENABLED";
    FD1S3AX multOut_i27 (.D(multOut_28__N_1217[27]), .CK(clk_N_683), .Q(multOut[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i27.GSR = "ENABLED";
    FD1S3AX multOut_i28 (.D(multOut_28__N_1217[28]), .CK(clk_N_683), .Q(multOut[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i28.GSR = "ENABLED";
    LUT4 i14_4_lut (.A(speed_set_m1[13]), .B(speed_set_m1[1]), .C(speed_set_m1[12]), 
         .D(speed_set_m1[2]), .Z(n35_adj_2142)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(speed_set_m1[15]), .B(n38), .C(n32), .D(speed_set_m1[10]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut (.A(n9_adj_2143), .B(n7_adj_2144), .C(n1349[10]), .D(n1349[13]), 
         .Z(n30_adj_2145)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i3_2_lut (.A(n1349[14]), .B(n1349[12]), .Z(n9_adj_2143)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_54 (.A(n1349[11]), .B(n1349[9]), .C(n10_adj_2146), 
         .D(n1349[7]), .Z(n7_adj_2144)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_54.init = 16'haaa8;
    LUT4 i4_4_lut_adj_55 (.A(n1349[6]), .B(n8_adj_2147), .C(n1349[4]), 
         .D(n4_adj_2148), .Z(n10_adj_2146)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_55.init = 16'hfeee;
    LUT4 i2_2_lut_adj_56 (.A(n1349[5]), .B(n1349[8]), .Z(n8_adj_2147)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_56.init = 16'heeee;
    LUT4 i1_4_lut_adj_57 (.A(n1349[3]), .B(n1349[2]), .C(n1349[1]), .D(n1349[0]), 
         .Z(n4_adj_2148)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_57.init = 16'haaa8;
    LUT4 mux_237_i8_3_lut_4_lut_3_lut (.A(n30_adj_2140), .B(n1307[15]), 
         .C(n2261[7]), .Z(n1443[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[25:42])
    defparam mux_237_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_135_i25_4_lut (.A(backOut2[24]), .B(backOut3[24]), .C(n21321), 
         .D(n9), .Z(n551[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i25_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_58 (.A(n9_adj_2149), .B(n7_adj_2150), .C(n1328[10]), 
         .D(n1328[13]), .Z(n30_adj_2141)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_58.init = 16'h8000;
    LUT4 i3_2_lut_adj_59 (.A(n1328[14]), .B(n1328[12]), .Z(n9_adj_2149)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_59.init = 16'h8888;
    LUT4 i1_4_lut_adj_60 (.A(n1328[11]), .B(n1328[9]), .C(n10_adj_2151), 
         .D(n1328[7]), .Z(n7_adj_2150)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_60.init = 16'haaa8;
    LUT4 i4_4_lut_adj_61 (.A(n1328[6]), .B(n8_adj_2152), .C(n1328[4]), 
         .D(n4_adj_2153), .Z(n10_adj_2151)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_61.init = 16'hfeee;
    LUT4 i2_2_lut_adj_62 (.A(n1328[5]), .B(n1328[8]), .Z(n8_adj_2152)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_62.init = 16'heeee;
    LUT4 i1_4_lut_adj_63 (.A(n1328[3]), .B(n1328[2]), .C(n1328[1]), .D(n1328[0]), 
         .Z(n4_adj_2153)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_63.init = 16'haaa8;
    FD1P3AX Out0_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i1.GSR = "ENABLED";
    FD1P3AX Out0_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_98), .CK(clk_N_683), 
            .Q(Out0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i2.GSR = "ENABLED";
    FD1P3AX Out0_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i3.GSR = "ENABLED";
    FD1P3AX Out0_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i4.GSR = "ENABLED";
    FD1P3AX Out0_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i5.GSR = "ENABLED";
    FD1P3AX Out0_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i6.GSR = "ENABLED";
    FD1P3AX Out0_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i7.GSR = "ENABLED";
    FD1P3AX Out0_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i8.GSR = "ENABLED";
    FD1P3AX Out0_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i9.GSR = "ENABLED";
    FD1P3AX Out0_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i10.GSR = "ENABLED";
    FD1P3AX Out0_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i11.GSR = "ENABLED";
    FD1P3AX Out0_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i12.GSR = "ENABLED";
    FD1P3AX Out0_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i13.GSR = "ENABLED";
    FD1P3AX Out0_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i14.GSR = "ENABLED";
    FD1P3AX Out0_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i15.GSR = "ENABLED";
    FD1P3AX Out0_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i16.GSR = "ENABLED";
    FD1P3AX Out0_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i17.GSR = "ENABLED";
    FD1P3AX Out0_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i18.GSR = "ENABLED";
    FD1P3AX Out0_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i19.GSR = "ENABLED";
    FD1P3AX Out0_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i20.GSR = "ENABLED";
    FD1P3AX Out0_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i21.GSR = "ENABLED";
    FD1P3AX Out0_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i22.GSR = "ENABLED";
    FD1P3AX Out0_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i23.GSR = "ENABLED";
    FD1P3AX Out0_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i24.GSR = "ENABLED";
    FD1P3AX Out0_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i25.GSR = "ENABLED";
    FD1P3AX Out0_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i26.GSR = "ENABLED";
    FD1P3AX Out0_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i27.GSR = "ENABLED";
    FD1P3AX Out0_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_98), 
            .CK(clk_N_683), .Q(Out0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i28.GSR = "ENABLED";
    FD1P3AX Out1_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i1.GSR = "ENABLED";
    FD1P3AX Out1_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_126), .CK(clk_N_683), 
            .Q(Out1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i2.GSR = "ENABLED";
    FD1P3AX Out1_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i3.GSR = "ENABLED";
    FD1P3AX Out1_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i4.GSR = "ENABLED";
    FD1P3AX Out1_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i5.GSR = "ENABLED";
    FD1P3AX Out1_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i6.GSR = "ENABLED";
    FD1P3AX Out1_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i7.GSR = "ENABLED";
    FD1P3AX Out1_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i8.GSR = "ENABLED";
    FD1P3AX Out1_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i9.GSR = "ENABLED";
    FD1P3AX Out1_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i10.GSR = "ENABLED";
    FD1P3AX Out1_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i11.GSR = "ENABLED";
    FD1P3AX Out1_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i12.GSR = "ENABLED";
    FD1P3AX Out1_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i13.GSR = "ENABLED";
    FD1P3AX Out1_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i14.GSR = "ENABLED";
    FD1P3AX Out1_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i15.GSR = "ENABLED";
    FD1P3AX Out1_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i16.GSR = "ENABLED";
    FD1P3AX Out1_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i17.GSR = "ENABLED";
    FD1P3AX Out1_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i18.GSR = "ENABLED";
    FD1P3AX Out1_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i19.GSR = "ENABLED";
    FD1P3AX Out1_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i20.GSR = "ENABLED";
    FD1P3AX Out1_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i21.GSR = "ENABLED";
    FD1P3AX Out1_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i22.GSR = "ENABLED";
    FD1P3AX Out1_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i23.GSR = "ENABLED";
    FD1P3AX Out1_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i24.GSR = "ENABLED";
    FD1P3AX Out1_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i25.GSR = "ENABLED";
    FD1P3AX Out1_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i26.GSR = "ENABLED";
    FD1P3AX Out1_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i27.GSR = "ENABLED";
    FD1P3AX Out1_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_126), 
            .CK(clk_N_683), .Q(Out1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i28.GSR = "ENABLED";
    FD1P3AX Out2_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i1.GSR = "ENABLED";
    FD1P3AX Out2_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_154), .CK(clk_N_683), 
            .Q(Out2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i2.GSR = "ENABLED";
    FD1P3AX Out2_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i3.GSR = "ENABLED";
    FD1P3AX Out2_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i4.GSR = "ENABLED";
    FD1P3AX Out2_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i5.GSR = "ENABLED";
    FD1P3AX Out2_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i6.GSR = "ENABLED";
    FD1P3AX Out2_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i7.GSR = "ENABLED";
    FD1P3AX Out2_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i8.GSR = "ENABLED";
    FD1P3AX Out2_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i9.GSR = "ENABLED";
    FD1P3AX Out2_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i10.GSR = "ENABLED";
    FD1P3AX Out2_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i11.GSR = "ENABLED";
    FD1P3AX Out2_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i12.GSR = "ENABLED";
    FD1P3AX Out2_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i13.GSR = "ENABLED";
    FD1P3AX Out2_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i14.GSR = "ENABLED";
    FD1P3AX Out2_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i15.GSR = "ENABLED";
    FD1P3AX Out2_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i16.GSR = "ENABLED";
    FD1P3AX Out2_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i17.GSR = "ENABLED";
    FD1P3AX Out2_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i18.GSR = "ENABLED";
    FD1P3AX Out2_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i19.GSR = "ENABLED";
    FD1P3AX Out2_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i20.GSR = "ENABLED";
    FD1P3AX Out2_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i21.GSR = "ENABLED";
    FD1P3AX Out2_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i22.GSR = "ENABLED";
    FD1P3AX Out2_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i23.GSR = "ENABLED";
    FD1P3AX Out2_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i24.GSR = "ENABLED";
    FD1P3AX Out2_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i25.GSR = "ENABLED";
    FD1P3AX Out2_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i26.GSR = "ENABLED";
    FD1P3AX Out2_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i27.GSR = "ENABLED";
    FD1P3AX Out2_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_154), 
            .CK(clk_N_683), .Q(Out2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i28.GSR = "ENABLED";
    FD1P3AX Out3_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i1.GSR = "ENABLED";
    FD1P3AX Out3_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_182), .CK(clk_N_683), 
            .Q(Out3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i2.GSR = "ENABLED";
    FD1P3AX Out3_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i3.GSR = "ENABLED";
    FD1P3AX Out3_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i4.GSR = "ENABLED";
    FD1P3AX Out3_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i5.GSR = "ENABLED";
    FD1P3AX Out3_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i6.GSR = "ENABLED";
    FD1P3AX Out3_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i7.GSR = "ENABLED";
    FD1P3AX Out3_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i8.GSR = "ENABLED";
    FD1P3AX Out3_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i9.GSR = "ENABLED";
    FD1P3AX Out3_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i10.GSR = "ENABLED";
    FD1P3AX Out3_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i11.GSR = "ENABLED";
    FD1P3AX Out3_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i12.GSR = "ENABLED";
    FD1P3AX Out3_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i13.GSR = "ENABLED";
    FD1P3AX Out3_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i14.GSR = "ENABLED";
    FD1P3AX Out3_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i15.GSR = "ENABLED";
    FD1P3AX Out3_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i16.GSR = "ENABLED";
    FD1P3AX Out3_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i17.GSR = "ENABLED";
    FD1P3AX Out3_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i18.GSR = "ENABLED";
    FD1P3AX Out3_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i19.GSR = "ENABLED";
    FD1P3AX Out3_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i20.GSR = "ENABLED";
    FD1P3AX Out3_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i21.GSR = "ENABLED";
    FD1P3AX Out3_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i22.GSR = "ENABLED";
    FD1P3AX Out3_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i23.GSR = "ENABLED";
    FD1P3AX Out3_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i24.GSR = "ENABLED";
    FD1P3AX Out3_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i25.GSR = "ENABLED";
    FD1P3AX Out3_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i26.GSR = "ENABLED";
    FD1P3AX Out3_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i27.GSR = "ENABLED";
    FD1P3AX Out3_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_182), 
            .CK(clk_N_683), .Q(Out3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i28.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_210), 
            .CK(clk_N_683), .Q(backOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i1 (.D(backOut3_28__N_1678[1]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i2 (.D(Out3_28__N_982[2]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i3 (.D(backOut3_28__N_1678[3]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i4 (.D(backOut3_28__N_1678[4]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i5 (.D(backOut3_28__N_1678[5]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i6 (.D(backOut3_28__N_1678[6]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i7 (.D(backOut3_28__N_1678[7]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i8 (.D(backOut3_28__N_1678[8]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i9 (.D(backOut3_28__N_1678[9]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i10 (.D(backOut3_28__N_1678[10]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i11 (.D(backOut3_28__N_1678[11]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i12 (.D(backOut3_28__N_1678[12]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i13 (.D(backOut3_28__N_1678[13]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i14 (.D(backOut3_28__N_1678[14]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i15 (.D(backOut3_28__N_1678[15]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i16 (.D(backOut3_28__N_1678[16]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i17 (.D(backOut3_28__N_1678[17]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i18 (.D(backOut3_28__N_1678[18]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i19 (.D(Out2_28__N_953[19]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i20 (.D(backOut3_28__N_1678[20]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i21 (.D(backOut3_28__N_1678[21]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i22 (.D(Out2_28__N_953[22]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i23 (.D(backOut3_28__N_1678[23]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i24 (.D(Out2_28__N_953[24]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i25 (.D(Out2_28__N_953[25]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i26 (.D(backOut3_28__N_1678[26]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i27 (.D(backOut3_28__N_1678[27]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i28 (.D(backOut2_28__N_1649[28]), .SP(clk_N_683_enable_238), 
            .CK(clk_N_683), .Q(backOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i28.GSR = "DISABLED";
    LUT4 i5_4_lut_adj_64 (.A(n9_adj_2154), .B(n7_adj_2155), .C(n1307[10]), 
         .D(n1307[13]), .Z(n30_adj_2140)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_64.init = 16'h8000;
    LUT4 i3_2_lut_adj_65 (.A(n1307[14]), .B(n1307[12]), .Z(n9_adj_2154)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_65.init = 16'h8888;
    LUT4 i1_4_lut_adj_66 (.A(n1307[11]), .B(n1307[9]), .C(n10_adj_2156), 
         .D(n1307[7]), .Z(n7_adj_2155)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_66.init = 16'haaa8;
    LUT4 i4_4_lut_adj_67 (.A(n1307[6]), .B(n8_adj_2157), .C(n1307[4]), 
         .D(n4_adj_2158), .Z(n10_adj_2156)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_67.init = 16'hfeee;
    LUT4 i2_2_lut_adj_68 (.A(n1307[5]), .B(n1307[8]), .Z(n8_adj_2157)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_68.init = 16'heeee;
    LUT4 i1_4_lut_adj_69 (.A(n1307[3]), .B(n1307[2]), .C(n1307[1]), .D(n1307[0]), 
         .Z(n4_adj_2158)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_69.init = 16'haaa8;
    LUT4 mux_135_i26_4_lut (.A(backOut2[25]), .B(backOut3[25]), .C(n21321), 
         .D(n9), .Z(n551[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i26_4_lut.init = 16'h0aca;
    FD1S3AX subOut_i1 (.D(\subOut_24__N_1177[1] ), .CK(clk_N_683), .Q(subOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i1.GSR = "ENABLED";
    FD1S3AX subOut_i2 (.D(\subOut_24__N_1177[2] ), .CK(clk_N_683), .Q(subOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i2.GSR = "ENABLED";
    FD1S3AX subOut_i3 (.D(\subOut_24__N_1177[3] ), .CK(clk_N_683), .Q(subOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i3.GSR = "ENABLED";
    FD1S3AX subOut_i4 (.D(\subOut_24__N_1177[4] ), .CK(clk_N_683), .Q(subOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i4.GSR = "ENABLED";
    FD1S3AX subOut_i5 (.D(\subOut_24__N_1177[5] ), .CK(clk_N_683), .Q(subOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i5.GSR = "ENABLED";
    FD1S3AX subOut_i6 (.D(\subOut_24__N_1177[6] ), .CK(clk_N_683), .Q(subOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i6.GSR = "ENABLED";
    FD1S3AX subOut_i7 (.D(\subOut_24__N_1177[7] ), .CK(clk_N_683), .Q(subOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i7.GSR = "ENABLED";
    FD1S3AX subOut_i8 (.D(\subOut_24__N_1177[8] ), .CK(clk_N_683), .Q(subOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i8.GSR = "ENABLED";
    FD1S3AX subOut_i9 (.D(\subOut_24__N_1177[9] ), .CK(clk_N_683), .Q(subOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i9.GSR = "ENABLED";
    FD1S3AX subOut_i10 (.D(\subOut_24__N_1177[10] ), .CK(clk_N_683), .Q(subOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i10.GSR = "ENABLED";
    FD1S3AX subOut_i11 (.D(\subOut_24__N_1177[11] ), .CK(clk_N_683), .Q(subOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i11.GSR = "ENABLED";
    FD1S3AX subOut_i12 (.D(\subOut_24__N_1177[12] ), .CK(clk_N_683), .Q(subOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i12.GSR = "ENABLED";
    FD1S3AX subOut_i13 (.D(\subOut_24__N_1177[13] ), .CK(clk_N_683), .Q(subOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i13.GSR = "ENABLED";
    FD1S3AX subOut_i14 (.D(\subOut_24__N_1177[14] ), .CK(clk_N_683), .Q(subOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i14.GSR = "ENABLED";
    FD1S3AX subOut_i15 (.D(\subOut_24__N_1177[15] ), .CK(clk_N_683), .Q(subOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i15.GSR = "ENABLED";
    FD1S3AX subOut_i16 (.D(\subOut_24__N_1177[16] ), .CK(clk_N_683), .Q(subOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i16.GSR = "ENABLED";
    FD1S3AX subOut_i17 (.D(\subOut_24__N_1177[17] ), .CK(clk_N_683), .Q(subOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i17.GSR = "ENABLED";
    FD1S3AX subOut_i18 (.D(\subOut_24__N_1177[18] ), .CK(clk_N_683), .Q(subOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i18.GSR = "ENABLED";
    FD1S3AX subOut_i19 (.D(\subOut_24__N_1177[19] ), .CK(clk_N_683), .Q(subOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i19.GSR = "ENABLED";
    FD1S3AX subOut_i20 (.D(\subOut_24__N_1177[20] ), .CK(clk_N_683), .Q(subOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i20.GSR = "ENABLED";
    FD1S3AX subOut_i21 (.D(\subOut_24__N_1177[21] ), .CK(clk_N_683), .Q(subOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i21.GSR = "ENABLED";
    FD1S3AX subOut_i23 (.D(\subOut_24__N_1177[24] ), .CK(clk_N_683), .Q(subOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i23.GSR = "ENABLED";
    LUT4 i5_4_lut_adj_70 (.A(n9_adj_2159), .B(n7_adj_2160), .C(n1286[10]), 
         .D(n1286[13]), .Z(n30)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_70.init = 16'h8000;
    LUT4 i3_2_lut_adj_71 (.A(n1286[14]), .B(n1286[12]), .Z(n9_adj_2159)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_71.init = 16'h8888;
    LUT4 i1_4_lut_adj_72 (.A(n1286[11]), .B(n1286[9]), .C(n10_adj_2161), 
         .D(n1286[7]), .Z(n7_adj_2160)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_72.init = 16'haaa8;
    LUT4 i4_4_lut_adj_73 (.A(n1286[6]), .B(n8_adj_2162), .C(n1286[4]), 
         .D(n4_adj_2163), .Z(n10_adj_2161)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_73.init = 16'hfeee;
    LUT4 i2_2_lut_adj_74 (.A(n1286[5]), .B(n1286[8]), .Z(n8_adj_2162)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_74.init = 16'heeee;
    LUT4 i1_4_lut_adj_75 (.A(n1286[3]), .B(n1286[2]), .C(n1286[1]), .D(n1286[0]), 
         .Z(n4_adj_2163)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_75.init = 16'haaa8;
    LUT4 i1_4_lut_adj_76 (.A(ss[3]), .B(n19508), .C(n22105), .D(n11489), 
         .Z(clk_N_683_enable_42)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_76.init = 16'hc4c0;
    LUT4 i11782_3_lut_4_lut (.A(n1328[15]), .B(n30_adj_2141), .C(n16394), 
         .D(clk_N_683_enable_392), .Z(n14352)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(362[7:42])
    defparam i11782_3_lut_4_lut.init = 16'hf700;
    LUT4 mux_135_i27_4_lut (.A(backOut2[26]), .B(backOut3[26]), .C(n21321), 
         .D(n9), .Z(n551[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i27_4_lut.init = 16'h0aca;
    LUT4 i15_4_lut (.A(speed_set_m1[0]), .B(speed_set_m1[7]), .C(speed_set_m1[17]), 
         .D(speed_set_m1[11]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i1816_1_lut (.A(ss[0]), .Z(n1)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1816_1_lut.init = 16'h5555;
    LUT4 mux_244_i7_3_lut_4_lut_3_lut (.A(n30_adj_2141), .B(n1328[15]), 
         .C(n2273[6]), .Z(n1487[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(362[25:42])
    defparam mux_244_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 mux_135_i28_4_lut (.A(backOut2[27]), .B(backOut3[27]), .C(n21321), 
         .D(n9), .Z(n551[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i28_4_lut.init = 16'h0aca;
    LUT4 mux_244_i8_3_lut_4_lut_3_lut (.A(n30_adj_2141), .B(n1328[15]), 
         .C(n2273[7]), .Z(n1487[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(362[25:42])
    defparam mux_244_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i1_4_lut_adj_77 (.A(ss[3]), .B(n19508), .C(n22105), .D(n19513), 
         .Z(clk_N_683_enable_70)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_77.init = 16'hc4c0;
    LUT4 i13241_2_lut (.A(addOut[0]), .B(n22105), .Z(Out3_28__N_982[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13241_2_lut.init = 16'h2222;
    LUT4 i2_3_lut_4_lut (.A(ss[0]), .B(n21356), .C(ss[3]), .D(n22105), 
         .Z(n19420)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0080;
    LUT4 i11796_2_lut_4_lut (.A(ss[3]), .B(n21353), .C(ss[1]), .D(clk_N_683_enable_392), 
         .Z(n14338)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11796_2_lut_4_lut.init = 16'hfe00;
    LUT4 i3066_3_lut (.A(n3832), .B(n1061), .C(addOut[28]), .Z(intgOut0_28__N_1433[28])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3066_3_lut.init = 16'h3232;
    LUT4 i3072_3_lut (.A(n3832), .B(n1061), .C(addOut[27]), .Z(intgOut0_28__N_1433[27])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3072_3_lut.init = 16'h3232;
    LUT4 i3076_3_lut (.A(n3832), .B(n1061), .C(addOut[26]), .Z(intgOut0_28__N_1433[26])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3076_3_lut.init = 16'h3232;
    LUT4 i3080_3_lut (.A(n3832), .B(n1061), .C(addOut[25]), .Z(intgOut0_28__N_1433[25])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3080_3_lut.init = 16'h3232;
    LUT4 i3088_3_lut (.A(n3832), .B(n1061), .C(addOut[24]), .Z(intgOut0_28__N_1433[24])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3088_3_lut.init = 16'h3232;
    LUT4 i3094_3_lut (.A(n3832), .B(n1061), .C(addOut[23]), .Z(intgOut0_28__N_1433[23])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3094_3_lut.init = 16'h3232;
    LUT4 i3096_3_lut (.A(n3832), .B(n1061), .C(addOut[22]), .Z(intgOut0_28__N_1433[22])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3096_3_lut.init = 16'h3232;
    LUT4 i3098_3_lut (.A(n3832), .B(n1061), .C(addOut[21]), .Z(intgOut0_28__N_1433[21])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3098_3_lut.init = 16'h3232;
    LUT4 i7_4_lut_adj_78 (.A(Out2[3]), .B(n14_adj_2164), .C(n10_adj_2165), 
         .D(Out2[4]), .Z(n18568)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i7_4_lut_adj_78.init = 16'hfffe;
    LUT4 i3100_3_lut (.A(n3832), .B(n1061), .C(addOut[20]), .Z(intgOut0_28__N_1433[20])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3100_3_lut.init = 16'h3232;
    LUT4 i6_4_lut_adj_79 (.A(Out2[11]), .B(Out2[7]), .C(Out2[2]), .D(Out2[10]), 
         .Z(n14_adj_2164)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i6_4_lut_adj_79.init = 16'hfffe;
    LUT4 i2_2_lut_adj_80 (.A(Out2[9]), .B(Out2[1]), .Z(n10_adj_2165)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i2_2_lut_adj_80.init = 16'heeee;
    LUT4 i4_4_lut_adj_81 (.A(Out2[5]), .B(Out2[6]), .C(Out2[0]), .D(n6_adj_2166), 
         .Z(n18569)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i4_4_lut_adj_81.init = 16'hfffe;
    LUT4 i1_2_lut_adj_82 (.A(Out2[8]), .B(Out2[12]), .Z(n6_adj_2166)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i1_2_lut_adj_82.init = 16'heeee;
    LUT4 i7_4_lut_adj_83 (.A(Out1[3]), .B(n14_adj_2167), .C(n10_adj_2168), 
         .D(Out1[4]), .Z(n18505)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i7_4_lut_adj_83.init = 16'hfffe;
    LUT4 i6_4_lut_adj_84 (.A(Out1[11]), .B(Out1[7]), .C(Out1[2]), .D(Out1[10]), 
         .Z(n14_adj_2167)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i6_4_lut_adj_84.init = 16'hfffe;
    LUT4 i2_2_lut_adj_85 (.A(Out1[9]), .B(Out1[1]), .Z(n10_adj_2168)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i2_2_lut_adj_85.init = 16'heeee;
    LUT4 i3058_3_lut (.A(n3832), .B(n1061), .C(addOut[15]), .Z(intgOut0_28__N_1433[15])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3058_3_lut.init = 16'h3232;
    LUT4 i3060_3_lut (.A(n3832), .B(n1061), .C(addOut[13]), .Z(intgOut0_28__N_1433[13])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3060_3_lut.init = 16'h3232;
    LUT4 i3064_3_lut (.A(n3832), .B(n1061), .C(addOut[12]), .Z(intgOut0_28__N_1433[12])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3064_3_lut.init = 16'h3232;
    LUT4 i3070_3_lut (.A(n3832), .B(n1061), .C(addOut[11]), .Z(intgOut0_28__N_1433[11])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3070_3_lut.init = 16'h3232;
    LUT4 i3074_3_lut (.A(n3832), .B(n1061), .C(addOut[10]), .Z(intgOut0_28__N_1433[10])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3074_3_lut.init = 16'h3232;
    LUT4 i3086_3_lut (.A(n3832), .B(n1061), .C(addOut[8]), .Z(intgOut0_28__N_1433[8])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3086_3_lut.init = 16'h3232;
    LUT4 i3092_3_lut (.A(n3832), .B(n1061), .C(addOut[7]), .Z(intgOut0_28__N_1433[7])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3092_3_lut.init = 16'h3232;
    LUT4 i1_4_lut_adj_86 (.A(n16536), .B(n19534), .C(n21337), .D(n22105), 
         .Z(clk_N_683_enable_390)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;
    defparam i1_4_lut_adj_86.init = 16'hf5dd;
    LUT4 i1_4_lut_adj_87 (.A(n3648), .B(n35_adj_2169), .C(n40_adj_2170), 
         .D(n36_adj_2171), .Z(n4_adj_2136)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_87.init = 16'haaa8;
    LUT4 i14_4_lut_adj_88 (.A(speed_set_m2[13]), .B(speed_set_m2[1]), .C(speed_set_m2[12]), 
         .D(speed_set_m2[2]), .Z(n35_adj_2169)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_88.init = 16'hfffe;
    LUT4 i19_4_lut_adj_89 (.A(speed_set_m2[15]), .B(n38_adj_2172), .C(n32_adj_2173), 
         .D(speed_set_m2[10]), .Z(n40_adj_2170)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_89.init = 16'hfffe;
    CCU2D add_219_7 (.A0(Out2[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18051), 
          .COUT(n18052), .S0(n1328[5]), .S1(n1328[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_7.INIT0 = 16'h5aaa;
    defparam add_219_7.INIT1 = 16'h5aaa;
    defparam add_219_7.INJECT1_0 = "NO";
    defparam add_219_7.INJECT1_1 = "NO";
    LUT4 i15_4_lut_adj_90 (.A(speed_set_m2[0]), .B(speed_set_m2[7]), .C(speed_set_m2[17]), 
         .D(speed_set_m2[11]), .Z(n36_adj_2171)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_90.init = 16'hfffe;
    LUT4 i17_4_lut (.A(speed_set_m2[8]), .B(n34), .C(n24), .D(speed_set_m2[16]), 
         .Z(n38_adj_2172)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(speed_set_m2[6]), .B(speed_set_m2[3]), .C(speed_set_m2[14]), 
         .Z(n32_adj_2173)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(speed_set_m2[20]), .B(speed_set_m2[19]), .C(speed_set_m2[9]), 
         .D(speed_set_m2[4]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut_adj_91 (.A(speed_set_m2[18]), .B(speed_set_m2[5]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_91.init = 16'heeee;
    LUT4 mux_135_i29_4_lut (.A(backOut2[28]), .B(backOut3[28]), .C(n21321), 
         .D(n9), .Z(n551[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i29_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_92 (.A(n16544), .B(n18492), .C(n21337), .D(n22105), 
         .Z(clk_N_683_enable_303)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;
    defparam i1_4_lut_adj_92.init = 16'hf5dd;
    CCU2D sub_16_rep_3_add_2_11 (.A0(n2341[9]), .B0(n4380), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[10]), .B1(n4379), .C1(GND_net), .D1(GND_net), 
          .CIN(n18127), .COUT(n18128), .S0(n4427), .S1(n4426));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_11.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_11.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_93 (.A(n3744), .B(n35_adj_2174), .C(n40_adj_2175), 
         .D(n36_adj_2176), .Z(n4_adj_2135)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_93.init = 16'haaa8;
    LUT4 i14_4_lut_adj_94 (.A(speed_set_m4[13]), .B(speed_set_m4[1]), .C(speed_set_m4[12]), 
         .D(speed_set_m4[2]), .Z(n35_adj_2174)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_94.init = 16'hfffe;
    LUT4 i4_4_lut_adj_95 (.A(Out1[5]), .B(Out1[6]), .C(Out1[0]), .D(n6_adj_2177), 
         .Z(n18506)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i4_4_lut_adj_95.init = 16'hfffe;
    LUT4 i1_2_lut_adj_96 (.A(Out1[8]), .B(Out1[12]), .Z(n6_adj_2177)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i1_2_lut_adj_96.init = 16'heeee;
    CCU2D add_15003_13 (.A0(speed_set_m1[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18343), .COUT(n18344));
    defparam add_15003_13.INIT0 = 16'hf555;
    defparam add_15003_13.INIT1 = 16'hf555;
    defparam add_15003_13.INJECT1_0 = "NO";
    defparam add_15003_13.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_9 (.A0(n2341[7]), .B0(n4382), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[8]), .B1(n4381), .C1(GND_net), .D1(GND_net), 
          .CIN(n18126), .COUT(n18127), .S0(n4429), .S1(n4428));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_9.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_9.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_9.INJECT1_1 = "NO";
    LUT4 i19_4_lut_adj_97 (.A(speed_set_m4[15]), .B(n38_adj_2178), .C(n32_adj_2179), 
         .D(speed_set_m4[10]), .Z(n40_adj_2175)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_97.init = 16'hfffe;
    LUT4 i15_4_lut_adj_98 (.A(speed_set_m4[0]), .B(speed_set_m4[7]), .C(speed_set_m4[17]), 
         .D(speed_set_m4[11]), .Z(n36_adj_2176)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_98.init = 16'hfffe;
    CCU2D sub_16_rep_3_add_2_7 (.A0(n2341[5]), .B0(n4384), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[6]), .B1(n4383), .C1(GND_net), .D1(GND_net), 
          .CIN(n18125), .COUT(n18126), .S0(n4431), .S1(n4430));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_7.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_7.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_7.INJECT1_1 = "NO";
    LUT4 i17_4_lut_adj_99 (.A(speed_set_m4[8]), .B(n34_adj_2180), .C(n24_adj_2181), 
         .D(speed_set_m4[16]), .Z(n38_adj_2178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_99.init = 16'hfffe;
    LUT4 i11_3_lut_adj_100 (.A(speed_set_m4[6]), .B(speed_set_m4[3]), .C(speed_set_m4[14]), 
         .Z(n32_adj_2179)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_100.init = 16'hfefe;
    LUT4 i13_4_lut_adj_101 (.A(speed_set_m4[20]), .B(speed_set_m4[19]), 
         .C(speed_set_m4[9]), .D(speed_set_m4[4]), .Z(n34_adj_2180)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_101.init = 16'hfffe;
    LUT4 i3_2_lut_adj_102 (.A(speed_set_m4[18]), .B(speed_set_m4[5]), .Z(n24_adj_2181)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_102.init = 16'heeee;
    CCU2D sub_16_rep_3_add_2_5 (.A0(n2341[3]), .B0(n4386), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[4]), .B1(n4385), .C1(GND_net), .D1(GND_net), 
          .CIN(n18124), .COUT(n18125), .S0(n4433), .S1(n4432));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_5.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_5.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_5.INJECT1_1 = "NO";
    LUT4 i17137_2_lut_3_lut_4_lut (.A(n22084), .B(n21359), .C(n4328), 
         .D(ss[2]), .Z(n20284)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i17137_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i7_4_lut_adj_103 (.A(Out0[3]), .B(n14_adj_2182), .C(n10_adj_2183), 
         .D(Out0[4]), .Z(n18586)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i7_4_lut_adj_103.init = 16'hfffe;
    LUT4 i6_4_lut_adj_104 (.A(Out0[11]), .B(Out0[7]), .C(Out0[2]), .D(Out0[10]), 
         .Z(n14_adj_2182)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i6_4_lut_adj_104.init = 16'hfffe;
    CCU2D sub_16_rep_3_add_2_3 (.A0(n2341[1]), .B0(n4388), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[2]), .B1(n4387), .C1(GND_net), .D1(GND_net), 
          .CIN(n18123), .COUT(n18124), .S0(n4435), .S1(n4434));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_3.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_3.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_3.INJECT1_1 = "NO";
    LUT4 i2_2_lut_adj_105 (.A(Out0[9]), .B(Out0[1]), .Z(n10_adj_2183)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i2_2_lut_adj_105.init = 16'heeee;
    CCU2D add_219_5 (.A0(Out2[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18050), 
          .COUT(n18051), .S0(n1328[3]), .S1(n1328[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_5.INIT0 = 16'h5aaa;
    defparam add_219_5.INIT1 = 16'h5aaa;
    defparam add_219_5.INJECT1_0 = "NO";
    defparam add_219_5.INJECT1_1 = "NO";
    CCU2D add_15003_11 (.A0(speed_set_m1[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18342), .COUT(n18343));
    defparam add_15003_11.INIT0 = 16'hf555;
    defparam add_15003_11.INIT1 = 16'hf555;
    defparam add_15003_11.INJECT1_0 = "NO";
    defparam add_15003_11.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[0]), .B1(n4389), .C1(GND_net), .D1(GND_net), 
          .COUT(n18123), .S1(n4436));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_1.INIT0 = 16'h0000;
    defparam sub_16_rep_3_add_2_1.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_1.INJECT1_1 = "NO";
    LUT4 i4_4_lut_adj_106 (.A(Out0[5]), .B(Out0[6]), .C(Out0[0]), .D(n6_adj_2184), 
         .Z(n18587)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i4_4_lut_adj_106.init = 16'hfffe;
    CCU2D add_219_3 (.A0(Out2[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18049), 
          .COUT(n18050), .S0(n1328[1]), .S1(n1328[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_3.INIT0 = 16'h5aaa;
    defparam add_219_3.INIT1 = 16'h5aaa;
    defparam add_219_3.INJECT1_0 = "NO";
    defparam add_219_3.INJECT1_1 = "NO";
    CCU2D add_219_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[13]), .B1(n18568), .C1(n18569), .D1(Out2[28]), .COUT(n18049), 
          .S1(n1328[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_1.INIT0 = 16'hF000;
    defparam add_219_1.INIT1 = 16'h56aa;
    defparam add_219_1.INJECT1_0 = "NO";
    defparam add_219_1.INJECT1_1 = "NO";
    CCU2D add_215_17 (.A0(Out1[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18048), 
          .S0(n1307[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_17.INIT0 = 16'h5aaa;
    defparam add_215_17.INIT1 = 16'h0000;
    defparam add_215_17.INJECT1_0 = "NO";
    defparam add_215_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_107 (.A(Out0[8]), .B(Out0[12]), .Z(n6_adj_2184)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i1_2_lut_adj_107.init = 16'heeee;
    LUT4 i1_2_lut_rep_370 (.A(ss[0]), .B(ss[3]), .Z(n21351)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_370.init = 16'heeee;
    LUT4 i2_2_lut_rep_353_3_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n21334)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_2_lut_rep_353_3_lut.init = 16'hefef;
    LUT4 i13664_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), .D(ss[2]), 
         .Z(n16214)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13664_2_lut_3_lut_4_lut.init = 16'hfeff;
    CCU2D add_215_15 (.A0(Out1[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18047), 
          .COUT(n18048), .S0(n1307[13]), .S1(n1307[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_15.INIT0 = 16'h5aaa;
    defparam add_215_15.INIT1 = 16'h5aaa;
    defparam add_215_15.INJECT1_0 = "NO";
    defparam add_215_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_108 (.A(ss[0]), .B(ss[2]), .C(ss[1]), .Z(n11489)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut_adj_108.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_109 (.A(ss[0]), .B(ss[2]), .C(ss[1]), .Z(n19513)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut_adj_109.init = 16'h0808;
    LUT4 i1_2_lut_rep_372 (.A(ss[0]), .B(n22099), .Z(n21353)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_372.init = 16'heeee;
    CCU2D add_215_13 (.A0(Out1[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18046), 
          .COUT(n18047), .S0(n1307[11]), .S1(n1307[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_13.INIT0 = 16'h5aaa;
    defparam add_215_13.INIT1 = 16'h5aaa;
    defparam add_215_13.INJECT1_0 = "NO";
    defparam add_215_13.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_110 (.A(ss[0]), .B(n22099), .C(ss[1]), .D(ss[3]), 
         .Z(n18492)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_3_lut_4_lut_adj_110.init = 16'h1000;
    LUT4 i13662_2_lut_3_lut_4_lut (.A(ss[0]), .B(n22099), .C(ss[1]), .D(ss[3]), 
         .Z(n16212)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13662_2_lut_3_lut_4_lut.init = 16'hfeff;
    CCU2D add_15003_9 (.A0(speed_set_m1[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18341), .COUT(n18342));
    defparam add_15003_9.INIT0 = 16'hf555;
    defparam add_15003_9.INIT1 = 16'h0aaa;
    defparam add_15003_9.INJECT1_0 = "NO";
    defparam add_15003_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_352_3_lut (.A(ss[0]), .B(ss[2]), .C(ss[3]), .Z(n21333)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_352_3_lut.init = 16'hefef;
    CCU2D add_215_11 (.A0(Out1[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18045), 
          .COUT(n18046), .S0(n1307[9]), .S1(n1307[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_11.INIT0 = 16'h5aaa;
    defparam add_215_11.INIT1 = 16'h5aaa;
    defparam add_215_11.INJECT1_0 = "NO";
    defparam add_215_11.INJECT1_1 = "NO";
    CCU2D add_15003_7 (.A0(speed_set_m1[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18340), .COUT(n18341));
    defparam add_15003_7.INIT0 = 16'h0aaa;
    defparam add_15003_7.INIT1 = 16'hf555;
    defparam add_15003_7.INJECT1_0 = "NO";
    defparam add_15003_7.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_356_4_lut (.A(ss[0]), .B(n22099), .C(ss[1]), .D(ss[3]), 
         .Z(n21337)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_3_lut_rep_356_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_111 (.A(n16540), .B(n16212), .C(n21337), .D(n22105), 
         .Z(clk_N_683_enable_331)) /* synthesis lut_function=((B (C (D))+!B (C+!(D)))+!A) */ ;
    defparam i1_4_lut_adj_111.init = 16'hf577;
    LUT4 i1_4_lut_adj_112 (.A(n3696), .B(n35_adj_2185), .C(n40_adj_2186), 
         .D(n36_adj_2187), .Z(n4)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_112.init = 16'haaa8;
    LUT4 i14_4_lut_adj_113 (.A(speed_set_m3[13]), .B(speed_set_m3[1]), .C(speed_set_m3[12]), 
         .D(speed_set_m3[2]), .Z(n35_adj_2185)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_113.init = 16'hfffe;
    CCU2D add_215_9 (.A0(Out1[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18044), 
          .COUT(n18045), .S0(n1307[7]), .S1(n1307[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_9.INIT0 = 16'h5aaa;
    defparam add_215_9.INIT1 = 16'h5aaa;
    defparam add_215_9.INJECT1_0 = "NO";
    defparam add_215_9.INJECT1_1 = "NO";
    LUT4 i19_4_lut_adj_114 (.A(speed_set_m3[15]), .B(n38_adj_2188), .C(n32_adj_2189), 
         .D(speed_set_m3[10]), .Z(n40_adj_2186)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_114.init = 16'hfffe;
    CCU2D add_215_7 (.A0(Out1[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18043), 
          .COUT(n18044), .S0(n1307[5]), .S1(n1307[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_7.INIT0 = 16'h5aaa;
    defparam add_215_7.INIT1 = 16'h5aaa;
    defparam add_215_7.INJECT1_0 = "NO";
    defparam add_215_7.INJECT1_1 = "NO";
    LUT4 i15_4_lut_adj_115 (.A(speed_set_m3[0]), .B(speed_set_m3[7]), .C(speed_set_m3[17]), 
         .D(speed_set_m3[11]), .Z(n36_adj_2187)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_115.init = 16'hfffe;
    LUT4 i17_4_lut_adj_116 (.A(speed_set_m3[8]), .B(n34_adj_2190), .C(n24_adj_2191), 
         .D(speed_set_m3[16]), .Z(n38_adj_2188)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_116.init = 16'hfffe;
    LUT4 i11_3_lut_adj_117 (.A(speed_set_m3[6]), .B(speed_set_m3[3]), .C(speed_set_m3[14]), 
         .Z(n32_adj_2189)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_117.init = 16'hfefe;
    CCU2D add_15003_5 (.A0(speed_set_m1[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18339), .COUT(n18340));
    defparam add_15003_5.INIT0 = 16'h0aaa;
    defparam add_15003_5.INIT1 = 16'h0aaa;
    defparam add_15003_5.INJECT1_0 = "NO";
    defparam add_15003_5.INJECT1_1 = "NO";
    LUT4 i13_4_lut_adj_118 (.A(speed_set_m3[20]), .B(speed_set_m3[19]), 
         .C(speed_set_m3[9]), .D(speed_set_m3[4]), .Z(n34_adj_2190)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_118.init = 16'hfffe;
    LUT4 i3_2_lut_adj_119 (.A(speed_set_m3[18]), .B(speed_set_m3[5]), .Z(n24_adj_2191)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_119.init = 16'heeee;
    LUT4 i11791_3_lut_4_lut (.A(n1349[15]), .B(n30_adj_2145), .C(n16394), 
         .D(clk_N_683_enable_392), .Z(n14361)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[7:42])
    defparam i11791_3_lut_4_lut.init = 16'hf700;
    LUT4 i3_4_lut (.A(n21294), .B(n21296), .C(n21295), .D(n16470), .Z(n11439)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i13351_2_lut (.A(addOut[5]), .B(n22105), .Z(backOut3_28__N_1678[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13351_2_lut.init = 16'h2222;
    LUT4 i2946_2_lut (.A(n22105), .B(n22100), .Z(clk_N_683_enable_392)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i2946_2_lut.init = 16'h8888;
    LUT4 i1743_1_lut (.A(n42), .Z(subIn1_24__N_1339)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(137[34:50])
    defparam i1743_1_lut.init = 16'h5555;
    LUT4 i1744_1_lut (.A(n49), .Z(dirout_m3_N_1753)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(139[35:51])
    defparam i1744_1_lut.init = 16'h5555;
    LUT4 i1742_1_lut (.A(n35), .Z(subIn1_24__N_1155)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(135[34:50])
    defparam i1742_1_lut.init = 16'h5555;
    LUT4 i13350_2_lut (.A(addOut[4]), .B(n22105), .Z(backOut3_28__N_1678[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13350_2_lut.init = 16'h2222;
    LUT4 i13349_2_lut (.A(addOut[3]), .B(n22105), .Z(backOut3_28__N_1678[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13349_2_lut.init = 16'h2222;
    CCU2D add_15003_3 (.A0(speed_set_m1[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18338), .COUT(n18339));
    defparam add_15003_3.INIT0 = 16'hf555;
    defparam add_15003_3.INIT1 = 16'hf555;
    defparam add_15003_3.INJECT1_0 = "NO";
    defparam add_15003_3.INJECT1_1 = "NO";
    CCU2D add_15003_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[4]), .B1(speed_set_m1[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18338));
    defparam add_15003_1.INIT0 = 16'hF000;
    defparam add_15003_1.INIT1 = 16'ha666;
    defparam add_15003_1.INJECT1_0 = "NO";
    defparam add_15003_1.INJECT1_1 = "NO";
    CCU2D add_15004_21 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18337), .S1(n49));
    defparam add_15004_21.INIT0 = 16'h5555;
    defparam add_15004_21.INIT1 = 16'h0000;
    defparam add_15004_21.INJECT1_0 = "NO";
    defparam add_15004_21.INJECT1_1 = "NO";
    CCU2D add_15004_19 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18336), .COUT(n18337));
    defparam add_15004_19.INIT0 = 16'hf555;
    defparam add_15004_19.INIT1 = 16'hf555;
    defparam add_15004_19.INJECT1_0 = "NO";
    defparam add_15004_19.INJECT1_1 = "NO";
    CCU2D add_215_5 (.A0(Out1[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18042), 
          .COUT(n18043), .S0(n1307[3]), .S1(n1307[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_5.INIT0 = 16'h5aaa;
    defparam add_215_5.INIT1 = 16'h5aaa;
    defparam add_215_5.INJECT1_0 = "NO";
    defparam add_215_5.INJECT1_1 = "NO";
    LUT4 i1745_1_lut (.A(n56), .Z(dirout_m4_N_1756)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(141[35:51])
    defparam i1745_1_lut.init = 16'h5555;
    CCU2D add_215_3 (.A0(Out1[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18041), 
          .COUT(n18042), .S0(n1307[1]), .S1(n1307[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_3.INIT0 = 16'h5aaa;
    defparam add_215_3.INIT1 = 16'h5aaa;
    defparam add_215_3.INJECT1_0 = "NO";
    defparam add_215_3.INJECT1_1 = "NO";
    LUT4 i13585_2_lut (.A(addOut[2]), .B(n22105), .Z(Out3_28__N_982[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13585_2_lut.init = 16'h2222;
    CCU2D add_215_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[13]), .B1(n18505), .C1(n18506), .D1(Out1[28]), .COUT(n18041), 
          .S1(n1307[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_1.INIT0 = 16'hF000;
    defparam add_215_1.INIT1 = 16'h56aa;
    defparam add_215_1.INJECT1_0 = "NO";
    defparam add_215_1.INJECT1_1 = "NO";
    CCU2D add_15004_17 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18335), .COUT(n18336));
    defparam add_15004_17.INIT0 = 16'hf555;
    defparam add_15004_17.INIT1 = 16'hf555;
    defparam add_15004_17.INJECT1_0 = "NO";
    defparam add_15004_17.INJECT1_1 = "NO";
    CCU2D add_211_17 (.A0(Out0[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18040), 
          .S0(n1286[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_17.INIT0 = 16'h5aaa;
    defparam add_211_17.INIT1 = 16'h0000;
    defparam add_211_17.INJECT1_0 = "NO";
    defparam add_211_17.INJECT1_1 = "NO";
    CCU2D add_211_15 (.A0(Out0[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18039), 
          .COUT(n18040), .S0(n1286[13]), .S1(n1286[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_15.INIT0 = 16'h5aaa;
    defparam add_211_15.INIT1 = 16'h5aaa;
    defparam add_211_15.INJECT1_0 = "NO";
    defparam add_211_15.INJECT1_1 = "NO";
    CCU2D add_211_13 (.A0(Out0[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18038), 
          .COUT(n18039), .S0(n1286[11]), .S1(n1286[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_13.INIT0 = 16'h5aaa;
    defparam add_211_13.INIT1 = 16'h5aaa;
    defparam add_211_13.INJECT1_0 = "NO";
    defparam add_211_13.INJECT1_1 = "NO";
    CCU2D add_15004_15 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18334), .COUT(n18335));
    defparam add_15004_15.INIT0 = 16'hf555;
    defparam add_15004_15.INIT1 = 16'hf555;
    defparam add_15004_15.INJECT1_0 = "NO";
    defparam add_15004_15.INJECT1_1 = "NO";
    CCU2D add_15004_13 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18333), .COUT(n18334));
    defparam add_15004_13.INIT0 = 16'hf555;
    defparam add_15004_13.INIT1 = 16'hf555;
    defparam add_15004_13.INJECT1_0 = "NO";
    defparam add_15004_13.INJECT1_1 = "NO";
    CCU2D add_15004_11 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18332), .COUT(n18333));
    defparam add_15004_11.INIT0 = 16'hf555;
    defparam add_15004_11.INIT1 = 16'hf555;
    defparam add_15004_11.INJECT1_0 = "NO";
    defparam add_15004_11.INJECT1_1 = "NO";
    CCU2D add_15004_9 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18331), .COUT(n18332));
    defparam add_15004_9.INIT0 = 16'hf555;
    defparam add_15004_9.INIT1 = 16'hf555;
    defparam add_15004_9.INJECT1_0 = "NO";
    defparam add_15004_9.INJECT1_1 = "NO";
    CCU2D add_211_11 (.A0(Out0[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18037), 
          .COUT(n18038), .S0(n1286[9]), .S1(n1286[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_11.INIT0 = 16'h5aaa;
    defparam add_211_11.INIT1 = 16'h5aaa;
    defparam add_211_11.INJECT1_0 = "NO";
    defparam add_211_11.INJECT1_1 = "NO";
    CCU2D add_211_9 (.A0(Out0[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18036), 
          .COUT(n18037), .S0(n1286[7]), .S1(n1286[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_9.INIT0 = 16'h5aaa;
    defparam add_211_9.INIT1 = 16'h5aaa;
    defparam add_211_9.INJECT1_0 = "NO";
    defparam add_211_9.INJECT1_1 = "NO";
    CCU2D add_15004_7 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18330), .COUT(n18331));
    defparam add_15004_7.INIT0 = 16'hf555;
    defparam add_15004_7.INIT1 = 16'hf555;
    defparam add_15004_7.INJECT1_0 = "NO";
    defparam add_15004_7.INJECT1_1 = "NO";
    CCU2D add_15004_5 (.A0(speed_set_m3[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18329), .COUT(n18330));
    defparam add_15004_5.INIT0 = 16'hf555;
    defparam add_15004_5.INIT1 = 16'hf555;
    defparam add_15004_5.INJECT1_0 = "NO";
    defparam add_15004_5.INJECT1_1 = "NO";
    CCU2D add_15004_3 (.A0(speed_set_m3[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18328), .COUT(n18329));
    defparam add_15004_3.INIT0 = 16'hf555;
    defparam add_15004_3.INIT1 = 16'hf555;
    defparam add_15004_3.INJECT1_0 = "NO";
    defparam add_15004_3.INJECT1_1 = "NO";
    CCU2D add_15004_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[0]), .B1(speed_set_m3[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18328));
    defparam add_15004_1.INIT0 = 16'hF000;
    defparam add_15004_1.INIT1 = 16'ha666;
    defparam add_15004_1.INJECT1_0 = "NO";
    defparam add_15004_1.INJECT1_1 = "NO";
    CCU2D add_15013_21 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18253), .S1(n56));
    defparam add_15013_21.INIT0 = 16'h5555;
    defparam add_15013_21.INIT1 = 16'h0000;
    defparam add_15013_21.INJECT1_0 = "NO";
    defparam add_15013_21.INJECT1_1 = "NO";
    LUT4 i13339_2_lut (.A(addOut[28]), .B(n22105), .Z(backOut2_28__N_1649[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13339_2_lut.init = 16'h2222;
    LUT4 i13409_2_lut (.A(addOut[27]), .B(n22105), .Z(backOut3_28__N_1678[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13409_2_lut.init = 16'h2222;
    CCU2D add_15013_19 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18252), .COUT(n18253));
    defparam add_15013_19.INIT0 = 16'hf555;
    defparam add_15013_19.INIT1 = 16'hf555;
    defparam add_15013_19.INJECT1_0 = "NO";
    defparam add_15013_19.INJECT1_1 = "NO";
    CCU2D add_15005_21 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18327), .S1(n42));
    defparam add_15005_21.INIT0 = 16'h5555;
    defparam add_15005_21.INIT1 = 16'h0000;
    defparam add_15005_21.INJECT1_0 = "NO";
    defparam add_15005_21.INJECT1_1 = "NO";
    CCU2D add_15005_19 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18326), .COUT(n18327));
    defparam add_15005_19.INIT0 = 16'hf555;
    defparam add_15005_19.INIT1 = 16'hf555;
    defparam add_15005_19.INJECT1_0 = "NO";
    defparam add_15005_19.INJECT1_1 = "NO";
    CCU2D add_15013_17 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18251), .COUT(n18252));
    defparam add_15013_17.INIT0 = 16'hf555;
    defparam add_15013_17.INIT1 = 16'hf555;
    defparam add_15013_17.INJECT1_0 = "NO";
    defparam add_15013_17.INJECT1_1 = "NO";
    CCU2D add_15005_17 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18325), .COUT(n18326));
    defparam add_15005_17.INIT0 = 16'hf555;
    defparam add_15005_17.INIT1 = 16'hf555;
    defparam add_15005_17.INJECT1_0 = "NO";
    defparam add_15005_17.INJECT1_1 = "NO";
    CCU2D add_15013_15 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18250), .COUT(n18251));
    defparam add_15013_15.INIT0 = 16'hf555;
    defparam add_15013_15.INIT1 = 16'hf555;
    defparam add_15013_15.INJECT1_0 = "NO";
    defparam add_15013_15.INJECT1_1 = "NO";
    CCU2D add_15013_13 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18249), .COUT(n18250));
    defparam add_15013_13.INIT0 = 16'hf555;
    defparam add_15013_13.INIT1 = 16'hf555;
    defparam add_15013_13.INJECT1_0 = "NO";
    defparam add_15013_13.INJECT1_1 = "NO";
    CCU2D add_211_7 (.A0(Out0[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18035), 
          .COUT(n18036), .S0(n1286[5]), .S1(n1286[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_7.INIT0 = 16'h5aaa;
    defparam add_211_7.INIT1 = 16'h5aaa;
    defparam add_211_7.INJECT1_0 = "NO";
    defparam add_211_7.INJECT1_1 = "NO";
    CCU2D add_15013_11 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18248), .COUT(n18249));
    defparam add_15013_11.INIT0 = 16'hf555;
    defparam add_15013_11.INIT1 = 16'hf555;
    defparam add_15013_11.INJECT1_0 = "NO";
    defparam add_15013_11.INJECT1_1 = "NO";
    CCU2D add_211_5 (.A0(Out0[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18034), 
          .COUT(n18035), .S0(n1286[3]), .S1(n1286[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_5.INIT0 = 16'h5aaa;
    defparam add_211_5.INIT1 = 16'h5aaa;
    defparam add_211_5.INJECT1_0 = "NO";
    defparam add_211_5.INJECT1_1 = "NO";
    CCU2D add_211_3 (.A0(Out0[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18033), 
          .COUT(n18034), .S0(n1286[1]), .S1(n1286[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_3.INIT0 = 16'h5aaa;
    defparam add_211_3.INIT1 = 16'h5aaa;
    defparam add_211_3.INJECT1_0 = "NO";
    defparam add_211_3.INJECT1_1 = "NO";
    CCU2D add_15005_15 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18324), .COUT(n18325));
    defparam add_15005_15.INIT0 = 16'hf555;
    defparam add_15005_15.INIT1 = 16'hf555;
    defparam add_15005_15.INJECT1_0 = "NO";
    defparam add_15005_15.INJECT1_1 = "NO";
    CCU2D add_15005_13 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18323), .COUT(n18324));
    defparam add_15005_13.INIT0 = 16'hf555;
    defparam add_15005_13.INIT1 = 16'hf555;
    defparam add_15005_13.INJECT1_0 = "NO";
    defparam add_15005_13.INJECT1_1 = "NO";
    CCU2D add_15013_9 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18247), .COUT(n18248));
    defparam add_15013_9.INIT0 = 16'hf555;
    defparam add_15013_9.INIT1 = 16'hf555;
    defparam add_15013_9.INJECT1_0 = "NO";
    defparam add_15013_9.INJECT1_1 = "NO";
    CCU2D add_15005_11 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18322), .COUT(n18323));
    defparam add_15005_11.INIT0 = 16'hf555;
    defparam add_15005_11.INIT1 = 16'hf555;
    defparam add_15005_11.INJECT1_0 = "NO";
    defparam add_15005_11.INJECT1_1 = "NO";
    CCU2D add_15005_9 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18321), .COUT(n18322));
    defparam add_15005_9.INIT0 = 16'hf555;
    defparam add_15005_9.INIT1 = 16'hf555;
    defparam add_15005_9.INJECT1_0 = "NO";
    defparam add_15005_9.INJECT1_1 = "NO";
    CCU2D add_211_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[13]), .B1(n18586), .C1(n18587), .D1(Out0[28]), .COUT(n18033), 
          .S1(n1286[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_1.INIT0 = 16'hF000;
    defparam add_211_1.INIT1 = 16'h56aa;
    defparam add_211_1.INJECT1_0 = "NO";
    defparam add_211_1.INJECT1_1 = "NO";
    CCU2D add_15013_7 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18246), .COUT(n18247));
    defparam add_15013_7.INIT0 = 16'hf555;
    defparam add_15013_7.INIT1 = 16'hf555;
    defparam add_15013_7.INJECT1_0 = "NO";
    defparam add_15013_7.INJECT1_1 = "NO";
    CCU2D add_15013_5 (.A0(speed_set_m4[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18245), .COUT(n18246));
    defparam add_15013_5.INIT0 = 16'hf555;
    defparam add_15013_5.INIT1 = 16'hf555;
    defparam add_15013_5.INJECT1_0 = "NO";
    defparam add_15013_5.INJECT1_1 = "NO";
    LUT4 i13347_2_lut (.A(addOut[1]), .B(n22105), .Z(backOut3_28__N_1678[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13347_2_lut.init = 16'h2222;
    CCU2D add_1176_23 (.A0(n5410), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18032), 
          .S0(n2341[21]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_23.INIT0 = 16'hf555;
    defparam add_1176_23.INIT1 = 16'h0000;
    defparam add_1176_23.INJECT1_0 = "NO";
    defparam add_1176_23.INJECT1_1 = "NO";
    FD1P3IX intgOut2_i0 (.D(addOut[0]), .SP(clk_N_683_enable_331), .CD(n14278), 
            .CK(clk_N_683), .Q(intgOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i0.GSR = "ENABLED";
    LUT4 i17_4_lut_adj_120 (.A(speed_set_m1[8]), .B(n34_adj_2192), .C(n24_adj_2193), 
         .D(speed_set_m1[16]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i17_4_lut_adj_120.init = 16'hfffe;
    LUT4 i11_3_lut_adj_121 (.A(speed_set_m1[6]), .B(speed_set_m1[3]), .C(speed_set_m1[14]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i11_3_lut_adj_121.init = 16'hfefe;
    CCU2D add_15005_7 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18320), .COUT(n18321));
    defparam add_15005_7.INIT0 = 16'hf555;
    defparam add_15005_7.INIT1 = 16'hf555;
    defparam add_15005_7.INJECT1_0 = "NO";
    defparam add_15005_7.INJECT1_1 = "NO";
    PFUMX mux_1190_i21 (.BLUT(n5362), .ALUT(n5320), .C0(n2533), .Z(n5410));
    PFUMX mux_1190_i20 (.BLUT(n5360), .ALUT(n5318), .C0(n2533), .Z(n5408));
    PFUMX mux_1190_i19 (.BLUT(n5358), .ALUT(n5316), .C0(n2533), .Z(n5406));
    PFUMX mux_1190_i18 (.BLUT(n5356), .ALUT(n5314), .C0(n2533), .Z(n5404));
    CCU2D add_15013_3 (.A0(speed_set_m4[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18244), .COUT(n18245));
    defparam add_15013_3.INIT0 = 16'hf555;
    defparam add_15013_3.INIT1 = 16'hf555;
    defparam add_15013_3.INJECT1_0 = "NO";
    defparam add_15013_3.INJECT1_1 = "NO";
    PFUMX mux_1190_i17 (.BLUT(n5354), .ALUT(n5312), .C0(n2533), .Z(n5402));
    PFUMX mux_1190_i16 (.BLUT(n5352), .ALUT(n5310), .C0(n2533), .Z(n5400));
    PFUMX mux_1190_i15 (.BLUT(n5350), .ALUT(n5308), .C0(n2533), .Z(n5398));
    PFUMX mux_1190_i14 (.BLUT(n5348), .ALUT(n5306), .C0(n2533), .Z(n5396));
    PFUMX mux_1190_i13 (.BLUT(n5346), .ALUT(n5304), .C0(n2533), .Z(n5394));
    PFUMX mux_1190_i12 (.BLUT(n5344), .ALUT(n5302), .C0(n2533), .Z(n5392));
    PFUMX mux_1190_i11 (.BLUT(n5342), .ALUT(n5300), .C0(n2533), .Z(n5390));
    PFUMX mux_1190_i10 (.BLUT(n5340), .ALUT(n5298), .C0(n2533), .Z(n5388));
    PFUMX mux_1190_i9 (.BLUT(n5338), .ALUT(n5296), .C0(n2533), .Z(n5386));
    CCU2D add_15005_5 (.A0(speed_set_m2[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18319), .COUT(n18320));
    defparam add_15005_5.INIT0 = 16'hf555;
    defparam add_15005_5.INIT1 = 16'hf555;
    defparam add_15005_5.INJECT1_0 = "NO";
    defparam add_15005_5.INJECT1_1 = "NO";
    PFUMX mux_1190_i8 (.BLUT(n5336), .ALUT(n5294), .C0(n2533), .Z(n5384));
    PFUMX mux_1190_i7 (.BLUT(n5334), .ALUT(n5292), .C0(n2533), .Z(n5382));
    PFUMX mux_1190_i6 (.BLUT(n5332), .ALUT(n5290), .C0(n2533), .Z(n5380));
    LUT4 i1_2_lut_rep_375 (.A(ss[1]), .B(ss[2]), .Z(n21356)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_375.init = 16'h8888;
    PFUMX mux_1190_i5 (.BLUT(n5330), .ALUT(n5288), .C0(n2533), .Z(n5378));
    LUT4 i9132_2_lut_3_lut_4_lut (.A(ss[1]), .B(ss[2]), .C(ss[3]), .D(ss[0]), 
         .Z(n15)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i9132_2_lut_3_lut_4_lut.init = 16'h78f0;
    PFUMX mux_1190_i4 (.BLUT(n5328), .ALUT(n5286), .C0(n2533), .Z(n5376));
    LUT4 i1_2_lut_3_lut_4_lut_adj_122 (.A(ss[1]), .B(n22099), .C(ss[3]), 
         .D(ss[0]), .Z(n19534)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_122.init = 16'h0008;
    PFUMX mux_1190_i3 (.BLUT(n5326), .ALUT(n5284), .C0(n2533), .Z(n5374));
    CCU2D add_15005_3 (.A0(speed_set_m2[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18318), .COUT(n18319));
    defparam add_15005_3.INIT0 = 16'hf555;
    defparam add_15005_3.INIT1 = 16'hf555;
    defparam add_15005_3.INJECT1_0 = "NO";
    defparam add_15005_3.INJECT1_1 = "NO";
    PFUMX mux_1190_i2 (.BLUT(n5324), .ALUT(n5282), .C0(n2533), .Z(n5372));
    CCU2D add_15005_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[0]), .B1(speed_set_m2[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18318));
    defparam add_15005_1.INIT0 = 16'hF000;
    defparam add_15005_1.INIT1 = 16'ha666;
    defparam add_15005_1.INJECT1_0 = "NO";
    defparam add_15005_1.INJECT1_1 = "NO";
    PFUMX mux_1190_i1 (.BLUT(n5280), .ALUT(n5278), .C0(n2533), .Z(n5370));
    PFUMX i3286 (.BLUT(n2581[1]), .ALUT(n5767), .C0(n21293), .Z(n5768));
    LUT4 i13406_2_lut (.A(addOut[26]), .B(n22105), .Z(backOut3_28__N_1678[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13406_2_lut.init = 16'h2222;
    PFUMX i3288 (.BLUT(n2581[2]), .ALUT(n5769), .C0(n21293), .Z(n5770));
    LUT4 i1815_2_lut_rep_378 (.A(ss[0]), .B(ss[1]), .Z(n21359)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1815_2_lut_rep_378.init = 16'h6666;
    PFUMX i3290 (.BLUT(n2581[3]), .ALUT(n5771), .C0(n21293), .Z(n5772));
    LUT4 i1_2_lut_rep_347_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n22099), 
         .D(n22084), .Z(n21328)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_347_3_lut_4_lut.init = 16'h0060;
    LUT4 i13578_2_lut (.A(addOut[25]), .B(n22105), .Z(Out2_28__N_953[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13578_2_lut.init = 16'h2222;
    PFUMX i3292 (.BLUT(n2581[4]), .ALUT(n5773), .C0(n21293), .Z(n5774));
    PFUMX i3294 (.BLUT(n2581[5]), .ALUT(n5775), .C0(n21293), .Z(n5776));
    PFUMX i3296 (.BLUT(n2581[6]), .ALUT(n5777), .C0(n21293), .Z(n5778));
    PFUMX i3298 (.BLUT(n2581[7]), .ALUT(n5779), .C0(n21293), .Z(n5780));
    CCU2D add_15013_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[0]), .B1(speed_set_m4[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18244));
    defparam add_15013_1.INIT0 = 16'hF000;
    defparam add_15013_1.INIT1 = 16'ha666;
    defparam add_15013_1.INJECT1_0 = "NO";
    defparam add_15013_1.INJECT1_1 = "NO";
    LUT4 i13577_2_lut (.A(addOut[24]), .B(n22105), .Z(Out2_28__N_953[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13577_2_lut.init = 16'h2222;
    PFUMX i3300 (.BLUT(n2581[8]), .ALUT(n5781), .C0(n21293), .Z(n5782));
    PFUMX i3302 (.BLUT(n2581[9]), .ALUT(n5783), .C0(n21293), .Z(n5784));
    PFUMX i3304 (.BLUT(n2581[10]), .ALUT(n5785), .C0(n21293), .Z(n5786));
    PFUMX i3306 (.BLUT(n2581[11]), .ALUT(n5787), .C0(n21293), .Z(n5788));
    PFUMX i3308 (.BLUT(n2581[12]), .ALUT(n5789), .C0(n21293), .Z(n5790));
    PFUMX i3310 (.BLUT(n2581[13]), .ALUT(n5791), .C0(n21293), .Z(n5792));
    PFUMX i3312 (.BLUT(n2581[14]), .ALUT(n5793), .C0(n21293), .Z(n5794));
    PFUMX i3314 (.BLUT(n2581[15]), .ALUT(n5795), .C0(n21293), .Z(n5796));
    PFUMX i3316 (.BLUT(n2581[16]), .ALUT(n5797), .C0(n21293), .Z(n5798));
    PFUMX i3318 (.BLUT(n2581[17]), .ALUT(n5799), .C0(n21293), .Z(n5800));
    PFUMX i3320 (.BLUT(n2581[18]), .ALUT(n5801), .C0(n21293), .Z(n5802));
    PFUMX i3322 (.BLUT(n2581[19]), .ALUT(n5803), .C0(n21293), .Z(n5804));
    PFUMX i3326 (.BLUT(n2581[20]), .ALUT(n5807), .C0(n21293), .Z(n5808));
    PFUMX i2999 (.BLUT(n2581[0]), .ALUT(n5480), .C0(n21293), .Z(n5481));
    L6MUX21 addIn2_28__I_29_i1 (.D0(n611[0]), .D1(addIn2_28__N_1375[0]), 
            .SD(n20045), .Z(addIn2_28__N_1246[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i2 (.D0(n611[1]), .D1(addIn2_28__N_1375[1]), 
            .SD(n20045), .Z(addIn2_28__N_1246[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i3 (.D0(n611[2]), .D1(addIn2_28__N_1375[2]), 
            .SD(n20045), .Z(addIn2_28__N_1246[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i4 (.D0(n611[3]), .D1(addIn2_28__N_1375[3]), 
            .SD(n20045), .Z(addIn2_28__N_1246[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i5 (.D0(n611[4]), .D1(addIn2_28__N_1375[4]), 
            .SD(n20045), .Z(addIn2_28__N_1246[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i6 (.D0(n611[5]), .D1(addIn2_28__N_1375[5]), 
            .SD(n20045), .Z(addIn2_28__N_1246[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i7 (.D0(n611[6]), .D1(addIn2_28__N_1375[6]), 
            .SD(n20045), .Z(addIn2_28__N_1246[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i8 (.D0(n611[7]), .D1(addIn2_28__N_1375[7]), 
            .SD(n20045), .Z(addIn2_28__N_1246[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i9 (.D0(n611[8]), .D1(addIn2_28__N_1375[8]), 
            .SD(n20045), .Z(addIn2_28__N_1246[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i10 (.D0(n611[9]), .D1(addIn2_28__N_1375[9]), 
            .SD(n20045), .Z(addIn2_28__N_1246[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i11 (.D0(n611[10]), .D1(addIn2_28__N_1375[10]), 
            .SD(n20045), .Z(addIn2_28__N_1246[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i12 (.D0(n611[11]), .D1(addIn2_28__N_1375[11]), 
            .SD(n20045), .Z(addIn2_28__N_1246[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i13 (.D0(n611[12]), .D1(addIn2_28__N_1375[12]), 
            .SD(n20045), .Z(addIn2_28__N_1246[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i14 (.D0(n611[13]), .D1(addIn2_28__N_1375[13]), 
            .SD(n20045), .Z(addIn2_28__N_1246[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i15 (.D0(n611[14]), .D1(addIn2_28__N_1375[14]), 
            .SD(n20045), .Z(addIn2_28__N_1246[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i16 (.D0(n611[15]), .D1(addIn2_28__N_1375[15]), 
            .SD(n20045), .Z(addIn2_28__N_1246[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13393_2_lut (.A(addOut[23]), .B(n22105), .Z(backOut3_28__N_1678[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13393_2_lut.init = 16'h2222;
    L6MUX21 addIn2_28__I_29_i17 (.D0(n611[16]), .D1(addIn2_28__N_1375[16]), 
            .SD(n20045), .Z(addIn2_28__N_1246[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i18 (.D0(n611[17]), .D1(addIn2_28__N_1375[17]), 
            .SD(n20045), .Z(addIn2_28__N_1246[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i19 (.D0(n611[18]), .D1(addIn2_28__N_1375[18]), 
            .SD(n20045), .Z(addIn2_28__N_1246[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i20 (.D0(n611[19]), .D1(addIn2_28__N_1375[19]), 
            .SD(n20045), .Z(addIn2_28__N_1246[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i21 (.D0(n611[20]), .D1(addIn2_28__N_1375[20]), 
            .SD(n20045), .Z(addIn2_28__N_1246[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i22 (.D0(n611[21]), .D1(addIn2_28__N_1375[21]), 
            .SD(n20045), .Z(addIn2_28__N_1246[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i23 (.D0(n611[22]), .D1(addIn2_28__N_1375[22]), 
            .SD(n20045), .Z(addIn2_28__N_1246[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i24 (.D0(n611[23]), .D1(addIn2_28__N_1375[23]), 
            .SD(n20045), .Z(addIn2_28__N_1246[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_251_i4_3_lut_4_lut_3_lut (.A(n30_adj_2145), .B(n1349[15]), 
         .C(n2285[3]), .Z(n1531[3])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[25:42])
    defparam mux_251_i4_3_lut_4_lut_3_lut.init = 16'hc4c4;
    L6MUX21 addIn2_28__I_29_i25 (.D0(n611[24]), .D1(addIn2_28__N_1375[24]), 
            .SD(n20045), .Z(addIn2_28__N_1246[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D sub_16_rep_4_add_2_23 (.A0(n8), .B0(n16260), .C0(n5808), .D0(n16270), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18243), 
          .S0(n4440));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_23.INIT0 = 16'h0f8f;
    defparam sub_16_rep_4_add_2_23.INIT1 = 16'h0000;
    defparam sub_16_rep_4_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_23.INJECT1_1 = "NO";
    L6MUX21 addIn2_28__I_29_i26 (.D0(n611[25]), .D1(addIn2_28__N_1375[25]), 
            .SD(n20045), .Z(addIn2_28__N_1246[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i27 (.D0(n611[26]), .D1(addIn2_28__N_1375[26]), 
            .SD(n20045), .Z(addIn2_28__N_1246[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i28 (.D0(n611[27]), .D1(addIn2_28__N_1375[27]), 
            .SD(n20045), .Z(addIn2_28__N_1246[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    L6MUX21 addIn2_28__I_29_i29 (.D0(n611[28]), .D1(addIn2_28__N_1375[28]), 
            .SD(n20045), .Z(addIn2_28__N_1246[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i19 (.BLUT(subIn2_24__N_1340[18]), .ALUT(subIn2_24__N_1156[18]), 
          .C0(n20284), .Z(n4371)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i18 (.BLUT(subIn2_24__N_1340[17]), .ALUT(subIn2_24__N_1156[17]), 
          .C0(n20284), .Z(n4372)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i17 (.BLUT(subIn2_24__N_1340[16]), .ALUT(subIn2_24__N_1156[16]), 
          .C0(n20284), .Z(n4373)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i16 (.BLUT(subIn2_24__N_1340[15]), .ALUT(subIn2_24__N_1156[15]), 
          .C0(n20284), .Z(n4374)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i15 (.BLUT(subIn2_24__N_1340[14]), .ALUT(subIn2_24__N_1156[14]), 
          .C0(n20284), .Z(n4375)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i14 (.BLUT(subIn2_24__N_1340[13]), .ALUT(subIn2_24__N_1156[13]), 
          .C0(n20284), .Z(n4376)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i13 (.BLUT(n367[12]), .ALUT(subIn2_24__N_1156[12]), 
          .C0(n20272), .Z(n4377)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i12 (.BLUT(subIn2_24__N_1340[11]), .ALUT(subIn2_24__N_1156[11]), 
          .C0(n20284), .Z(n4378)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13575_2_lut (.A(addOut[22]), .B(n22105), .Z(Out2_28__N_953[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13575_2_lut.init = 16'h2222;
    PFUMX subIn2_24__I_0_rep_1_i11 (.BLUT(subIn2_24__N_1340[10]), .ALUT(subIn2_24__N_1156[10]), 
          .C0(n20284), .Z(n4379)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D sub_16_rep_4_add_2_21 (.A0(n7), .B0(n11439), .C0(n5804), .D0(n16270), 
          .A1(n8), .B1(n16260), .C1(n5808), .D1(n16270), .CIN(n18242), 
          .COUT(n18243), .S0(n4442), .S1(n4441));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_21.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_21.INIT1 = 16'h0f8f;
    defparam sub_16_rep_4_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_21.INJECT1_1 = "NO";
    CCU2D add_15006_21 (.A0(speed_set_m1[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18317), .S1(n35));
    defparam add_15006_21.INIT0 = 16'h5555;
    defparam add_15006_21.INIT1 = 16'h0000;
    defparam add_15006_21.INJECT1_0 = "NO";
    defparam add_15006_21.INJECT1_1 = "NO";
    PFUMX subIn2_24__I_0_rep_1_i10 (.BLUT(n367[9]), .ALUT(subIn2_24__N_1156[9]), 
          .C0(n20272), .Z(n4380)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i9 (.BLUT(n367[8]), .ALUT(subIn2_24__N_1156[8]), 
          .C0(n20272), .Z(n4381)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i8 (.BLUT(n367[7]), .ALUT(subIn2_24__N_1156[7]), 
          .C0(n20272), .Z(n4382)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i7 (.BLUT(subIn2_24__N_1340[6]), .ALUT(subIn2_24__N_1156[6]), 
          .C0(n20284), .Z(n4383)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i6 (.BLUT(subIn2_24__N_1340[5]), .ALUT(subIn2_24__N_1156[5]), 
          .C0(n20284), .Z(n4384)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i5 (.BLUT(subIn2_24__N_1340[4]), .ALUT(subIn2_24__N_1156[4]), 
          .C0(n20284), .Z(n4385)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i4 (.BLUT(n367[3]), .ALUT(subIn2_24__N_1156[3]), 
          .C0(n20272), .Z(n4386)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i3 (.BLUT(subIn2_24__N_1340[2]), .ALUT(subIn2_24__N_1156[2]), 
          .C0(n20284), .Z(n4387)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i2 (.BLUT(subIn2_24__N_1340[1]), .ALUT(subIn2_24__N_1156[1]), 
          .C0(n20284), .Z(n4388)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX subIn2_24__I_0_rep_1_i1 (.BLUT(subIn2_24__N_1340[0]), .ALUT(subIn2_24__N_1156[0]), 
          .C0(n20284), .Z(n4389)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i2 (.BLUT(n551[1]), .ALUT(n671[1]), .C0(n20019), .Z(addIn2_28__N_1375[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i3 (.BLUT(n551[2]), .ALUT(n671[2]), .C0(n20019), .Z(addIn2_28__N_1375[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13385_2_lut (.A(addOut[21]), .B(n22105), .Z(backOut3_28__N_1678[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13385_2_lut.init = 16'h2222;
    LUT4 mux_251_i9_3_lut_4_lut_3_lut (.A(n30_adj_2145), .B(n1349[15]), 
         .C(n2285[8]), .Z(n1531[8])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[25:42])
    defparam mux_251_i9_3_lut_4_lut_3_lut.init = 16'hc4c4;
    PFUMX mux_140_i4 (.BLUT(n551[3]), .ALUT(n671[3]), .C0(n20019), .Z(addIn2_28__N_1375[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i5 (.BLUT(n551[4]), .ALUT(n671[4]), .C0(n20019), .Z(addIn2_28__N_1375[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i6 (.BLUT(n551[5]), .ALUT(n671[5]), .C0(n20019), .Z(addIn2_28__N_1375[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i7 (.BLUT(n551[6]), .ALUT(n671[6]), .C0(n20019), .Z(addIn2_28__N_1375[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i8 (.BLUT(n551[7]), .ALUT(n671[7]), .C0(n20019), .Z(addIn2_28__N_1375[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i9 (.BLUT(n551[8]), .ALUT(n671[8]), .C0(n20019), .Z(addIn2_28__N_1375[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i10 (.BLUT(n551[9]), .ALUT(n671[9]), .C0(n20019), .Z(addIn2_28__N_1375[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i11 (.BLUT(n551[10]), .ALUT(n671[10]), .C0(n20019), 
          .Z(addIn2_28__N_1375[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i12 (.BLUT(n551[11]), .ALUT(n671[11]), .C0(n20019), 
          .Z(addIn2_28__N_1375[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i13 (.BLUT(n551[12]), .ALUT(n671[12]), .C0(n20019), 
          .Z(addIn2_28__N_1375[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i14 (.BLUT(n551[13]), .ALUT(n671[13]), .C0(n20019), 
          .Z(addIn2_28__N_1375[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i15 (.BLUT(n551[14]), .ALUT(n671[14]), .C0(n20019), 
          .Z(addIn2_28__N_1375[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i16 (.BLUT(n551[15]), .ALUT(n671[15]), .C0(n20019), 
          .Z(addIn2_28__N_1375[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i17 (.BLUT(n551[16]), .ALUT(n671[16]), .C0(n20019), 
          .Z(addIn2_28__N_1375[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i18 (.BLUT(n551[17]), .ALUT(n671[17]), .C0(n20019), 
          .Z(addIn2_28__N_1375[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D sub_16_rep_4_add_2_19 (.A0(n4372), .B0(n11439), .C0(n5800), 
          .D0(n16270), .A1(n4371), .B1(n11439), .C1(n5802), .D1(n16270), 
          .CIN(n18241), .COUT(n18242), .S0(n4444), .S1(n4443));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_19.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_19.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_19.INJECT1_1 = "NO";
    PFUMX mux_140_i19 (.BLUT(n551[18]), .ALUT(n671[18]), .C0(n20019), 
          .Z(addIn2_28__N_1375[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i20 (.BLUT(n551[19]), .ALUT(n671[19]), .C0(n20019), 
          .Z(addIn2_28__N_1375[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13_4_lut_adj_123 (.A(speed_set_m1[20]), .B(speed_set_m1[19]), 
         .C(speed_set_m1[9]), .D(speed_set_m1[4]), .Z(n34_adj_2192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i13_4_lut_adj_123.init = 16'hfffe;
    CCU2D add_15006_19 (.A0(speed_set_m1[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18316), .COUT(n18317));
    defparam add_15006_19.INIT0 = 16'hf555;
    defparam add_15006_19.INIT1 = 16'hf555;
    defparam add_15006_19.INJECT1_0 = "NO";
    defparam add_15006_19.INJECT1_1 = "NO";
    PFUMX mux_140_i21 (.BLUT(n551[20]), .ALUT(n671[20]), .C0(n20019), 
          .Z(addIn2_28__N_1375[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i22 (.BLUT(n551[21]), .ALUT(n671[21]), .C0(n20019), 
          .Z(addIn2_28__N_1375[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_15006_17 (.A0(speed_set_m1[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18315), .COUT(n18316));
    defparam add_15006_17.INIT0 = 16'hf555;
    defparam add_15006_17.INIT1 = 16'hf555;
    defparam add_15006_17.INJECT1_0 = "NO";
    defparam add_15006_17.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_17 (.A0(n4374), .B0(n11439), .C0(n5796), 
          .D0(n16270), .A1(n4373), .B1(n11439), .C1(n5798), .D1(n16270), 
          .CIN(n18240), .COUT(n18241), .S0(n4446), .S1(n4445));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_17.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_17.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_17.INJECT1_1 = "NO";
    PFUMX mux_140_i1 (.BLUT(n551[0]), .ALUT(n671[0]), .C0(n20019), .Z(addIn2_28__N_1375[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13382_2_lut (.A(addOut[20]), .B(n22105), .Z(backOut3_28__N_1678[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13382_2_lut.init = 16'h2222;
    CCU2D add_15006_15 (.A0(speed_set_m1[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18314), .COUT(n18315));
    defparam add_15006_15.INIT0 = 16'hf555;
    defparam add_15006_15.INIT1 = 16'hf555;
    defparam add_15006_15.INJECT1_0 = "NO";
    defparam add_15006_15.INJECT1_1 = "NO";
    PFUMX mux_140_i23 (.BLUT(n551[22]), .ALUT(n671[22]), .C0(n20019), 
          .Z(addIn2_28__N_1375[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_140_i24 (.BLUT(n551[23]), .ALUT(n671[23]), .C0(n20019), 
          .Z(addIn2_28__N_1375[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX dutyout_m4_i0_i9 (.D(n1531[9]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i8 (.D(n1531[8]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i7 (.D(n1531[7]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i6 (.D(n1531[6]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i5 (.D(n1531[5]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i4 (.D(n2285[4]), .SP(clk_N_683_enable_392), .CD(n14361), 
            .CK(clk_N_683), .Q(PWMdut_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i3 (.D(n1531[3]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i3.GSR = "DISABLED";
    LUT4 i13572_2_lut (.A(addOut[19]), .B(n22105), .Z(Out2_28__N_953[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13572_2_lut.init = 16'h2222;
    PFUMX mux_140_i25 (.BLUT(n551[24]), .ALUT(n671[24]), .C0(n20019), 
          .Z(addIn2_28__N_1375[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX dutyout_m4_i0_i2 (.D(n2285[2]), .SP(clk_N_683_enable_392), .CD(n14361), 
            .CK(clk_N_683), .Q(PWMdut_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i1 (.D(n2285[1]), .SP(clk_N_683_enable_392), .CD(n14361), 
            .CK(clk_N_683), .Q(PWMdut_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i9 (.D(n1487[9]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i8 (.D(n1487[8]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i7 (.D(n1487[7]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i6 (.D(n1487[6]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i5 (.D(n1487[5]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i4 (.D(n2273[4]), .SP(clk_N_683_enable_392), .CD(n14352), 
            .CK(clk_N_683), .Q(PWMdut_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i3 (.D(n1487[3]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i2 (.D(n2273[2]), .SP(clk_N_683_enable_392), .CD(n14352), 
            .CK(clk_N_683), .Q(PWMdut_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i1 (.D(n2273[1]), .SP(clk_N_683_enable_392), .CD(n14352), 
            .CK(clk_N_683), .Q(PWMdut_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i9 (.D(n1443[9]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i9.GSR = "DISABLED";
    CCU2D sub_16_rep_4_add_2_15 (.A0(n4376), .B0(n11439), .C0(n5792), 
          .D0(n16270), .A1(n4375), .B1(n11439), .C1(n5794), .D1(n16270), 
          .CIN(n18239), .COUT(n18240), .S0(n4448), .S1(n4447));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_15.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_15.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_15.INJECT1_1 = "NO";
    FD1P3IX dutyout_m2_i0_i8 (.D(n1443[8]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i7 (.D(n1443[7]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i6 (.D(n1443[6]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i6.GSR = "DISABLED";
    PFUMX mux_140_i26 (.BLUT(n551[25]), .ALUT(n671[25]), .C0(n20019), 
          .Z(addIn2_28__N_1375[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX dutyout_m2_i0_i5 (.D(n1443[5]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i4 (.D(n2261[4]), .SP(clk_N_683_enable_392), .CD(n14343), 
            .CK(clk_N_683), .Q(PWMdut_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i3 (.D(n1443[3]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i3.GSR = "DISABLED";
    CCU2D sub_16_rep_4_add_2_13 (.A0(n4378), .B0(n11439), .C0(n5788), 
          .D0(n16270), .A1(n4377), .B1(n11439), .C1(n5790), .D1(n16270), 
          .CIN(n18238), .COUT(n18239), .S0(n4450), .S1(n4449));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_13.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_13.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_13.INJECT1_1 = "NO";
    FD1P3IX dutyout_m2_i0_i2 (.D(n2261[2]), .SP(clk_N_683_enable_392), .CD(n14343), 
            .CK(clk_N_683), .Q(PWMdut_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i1 (.D(n2261[1]), .SP(clk_N_683_enable_392), .CD(n14343), 
            .CK(clk_N_683), .Q(PWMdut_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i9 (.D(n1399[9]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i9.GSR = "DISABLED";
    PFUMX mux_140_i27 (.BLUT(n551[26]), .ALUT(n671[26]), .C0(n20019), 
          .Z(addIn2_28__N_1375[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX dutyout_m1_i0_i8 (.D(n1399[8]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i7 (.D(n1399[7]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i7.GSR = "DISABLED";
    CCU2D add_15006_13 (.A0(speed_set_m1[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18313), .COUT(n18314));
    defparam add_15006_13.INIT0 = 16'hf555;
    defparam add_15006_13.INIT1 = 16'hf555;
    defparam add_15006_13.INJECT1_0 = "NO";
    defparam add_15006_13.INJECT1_1 = "NO";
    FD1P3IX dutyout_m1_i0_i6 (.D(n1399[6]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i5 (.D(n1399[5]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i4 (.D(n2249[4]), .SP(clk_N_683_enable_392), .CD(n14334), 
            .CK(clk_N_683), .Q(PWMdut_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i3 (.D(n1399[3]), .SP(clk_N_683_enable_392), .CD(n14338), 
            .CK(clk_N_683), .Q(PWMdut_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i3.GSR = "DISABLED";
    LUT4 equal_133_i9_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21378), 
         .D(n22099), .Z(n9)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(164[29:36])
    defparam equal_133_i9_2_lut_3_lut_4_lut.init = 16'hfbff;
    PFUMX mux_140_i28 (.BLUT(n551[27]), .ALUT(n671[27]), .C0(n20019), 
          .Z(addIn2_28__N_1375[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX dutyout_m1_i0_i2 (.D(n2249[2]), .SP(clk_N_683_enable_392), .CD(n14334), 
            .CK(clk_N_683), .Q(PWMdut_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i1 (.D(n2249[1]), .SP(clk_N_683_enable_392), .CD(n14334), 
            .CK(clk_N_683), .Q(PWMdut_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i1.GSR = "DISABLED";
    FD1P3IX intgOut3_i28 (.D(intgOut0_28__N_1433[28]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i28.GSR = "ENABLED";
    FD1P3IX intgOut3_i27 (.D(intgOut0_28__N_1433[27]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i27.GSR = "ENABLED";
    FD1P3IX intgOut3_i26 (.D(intgOut0_28__N_1433[26]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i26.GSR = "ENABLED";
    FD1P3IX intgOut3_i25 (.D(intgOut0_28__N_1433[25]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i25.GSR = "ENABLED";
    FD1P3IX intgOut3_i24 (.D(intgOut0_28__N_1433[24]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i24.GSR = "ENABLED";
    LUT4 ss_4__I_0_358_i6_2_lut_rep_396 (.A(ss[0]), .B(ss[1]), .Z(n21377)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam ss_4__I_0_358_i6_2_lut_rep_396.init = 16'hdddd;
    FD1P3IX intgOut3_i23 (.D(intgOut0_28__N_1433[23]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i23.GSR = "ENABLED";
    FD1P3IX intgOut3_i22 (.D(intgOut0_28__N_1433[22]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i22.GSR = "ENABLED";
    FD1P3IX intgOut3_i21 (.D(intgOut0_28__N_1433[21]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i21.GSR = "ENABLED";
    FD1P3IX intgOut3_i20 (.D(intgOut0_28__N_1433[20]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i20.GSR = "ENABLED";
    FD1P3IX intgOut3_i19 (.D(intgOut0_28__N_1433[19]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i19.GSR = "ENABLED";
    FD1P3IX intgOut3_i18 (.D(intgOut0_28__N_1433[18]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i18.GSR = "ENABLED";
    FD1P3IX intgOut3_i17 (.D(intgOut0_28__N_1433[17]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i17.GSR = "ENABLED";
    FD1P3IX intgOut3_i16 (.D(intgOut0_28__N_1433[16]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i16.GSR = "ENABLED";
    LUT4 i17205_2_lut_rep_327_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21378), 
         .D(ss[2]), .Z(n21308)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam i17205_2_lut_rep_327_2_lut_3_lut_4_lut.init = 16'h0002;
    FD1P3IX intgOut3_i15 (.D(intgOut0_28__N_1433[15]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i15.GSR = "ENABLED";
    FD1P3IX intgOut3_i14 (.D(intgOut0_28__N_1433[14]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i14.GSR = "ENABLED";
    CCU2D sub_16_rep_4_add_2_11 (.A0(n4380), .B0(n11439), .C0(n5784), 
          .D0(n16270), .A1(n4379), .B1(n11439), .C1(n5786), .D1(n16270), 
          .CIN(n18237), .COUT(n18238), .S0(n4452), .S1(n4451));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_11.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_11.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_11.INJECT1_1 = "NO";
    FD1P3IX intgOut3_i13 (.D(intgOut0_28__N_1433[13]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i13.GSR = "ENABLED";
    FD1P3IX intgOut3_i12 (.D(intgOut0_28__N_1433[12]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i12.GSR = "ENABLED";
    FD1P3IX intgOut3_i11 (.D(intgOut0_28__N_1433[11]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i11.GSR = "ENABLED";
    FD1P3IX intgOut3_i10 (.D(intgOut0_28__N_1433[10]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i10.GSR = "ENABLED";
    FD1P3IX intgOut3_i9 (.D(intgOut0_28__N_1433[9]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i9.GSR = "ENABLED";
    FD1P3IX intgOut3_i8 (.D(intgOut0_28__N_1433[8]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i8.GSR = "ENABLED";
    FD1P3IX intgOut3_i7 (.D(intgOut0_28__N_1433[7]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i7.GSR = "ENABLED";
    LUT4 equal_114_i9_2_lut_rep_340_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21378), 
         .D(n22099), .Z(n21321)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam equal_114_i9_2_lut_rep_340_3_lut_4_lut.init = 16'hfdff;
    FD1P3IX intgOut3_i6 (.D(intgOut0_28__N_1433[6]), .SP(clk_N_683_enable_303), 
            .CD(n14312), .CK(clk_N_683), .Q(intgOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i6.GSR = "ENABLED";
    FD1P3IX intgOut3_i5 (.D(addOut[5]), .SP(clk_N_683_enable_303), .CD(n14307), 
            .CK(clk_N_683), .Q(intgOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i5.GSR = "ENABLED";
    FD1P3IX intgOut3_i4 (.D(addOut[4]), .SP(clk_N_683_enable_303), .CD(n14307), 
            .CK(clk_N_683), .Q(intgOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i4.GSR = "ENABLED";
    FD1P3IX intgOut3_i3 (.D(addOut[3]), .SP(clk_N_683_enable_303), .CD(n14307), 
            .CK(clk_N_683), .Q(intgOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i3.GSR = "ENABLED";
    FD1P3IX intgOut3_i2 (.D(addOut[2]), .SP(clk_N_683_enable_303), .CD(n14307), 
            .CK(clk_N_683), .Q(intgOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i2.GSR = "ENABLED";
    FD1P3IX intgOut3_i1 (.D(addOut[1]), .SP(clk_N_683_enable_303), .CD(n14307), 
            .CK(clk_N_683), .Q(intgOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i1.GSR = "ENABLED";
    FD1P3IX intgOut2_i28 (.D(intgOut0_28__N_1433[28]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i28.GSR = "ENABLED";
    FD1P3IX intgOut2_i27 (.D(intgOut0_28__N_1433[27]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i27.GSR = "ENABLED";
    FD1P3IX intgOut2_i26 (.D(intgOut0_28__N_1433[26]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i26.GSR = "ENABLED";
    LUT4 ss_4__I_0_358_i9_2_lut_rep_339_3_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n22084), .D(ss[2]), .Z(n21320)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam ss_4__I_0_358_i9_2_lut_rep_339_3_lut_4_lut.init = 16'hfdff;
    FD1P3IX intgOut2_i25 (.D(intgOut0_28__N_1433[25]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i25.GSR = "ENABLED";
    FD1P3IX intgOut2_i24 (.D(intgOut0_28__N_1433[24]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i24.GSR = "ENABLED";
    FD1P3IX intgOut2_i23 (.D(intgOut0_28__N_1433[23]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i23.GSR = "ENABLED";
    CCU2D sub_16_rep_4_add_2_9 (.A0(n4382), .B0(n11439), .C0(n5780), .D0(n16270), 
          .A1(n4381), .B1(n11439), .C1(n5782), .D1(n16270), .CIN(n18236), 
          .COUT(n18237), .S0(n4454), .S1(n4453));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_9.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_9.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_9.INJECT1_1 = "NO";
    FD1P3IX intgOut2_i22 (.D(intgOut0_28__N_1433[22]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i22.GSR = "ENABLED";
    FD1P3IX intgOut2_i21 (.D(intgOut0_28__N_1433[21]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i21.GSR = "ENABLED";
    FD1P3IX intgOut2_i20 (.D(intgOut0_28__N_1433[20]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i20.GSR = "ENABLED";
    CCU2D add_1176_21 (.A0(n5408), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5410), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18031), 
          .COUT(n18032), .S0(n2341[19]), .S1(n2341[20]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_21.INIT0 = 16'hf555;
    defparam add_1176_21.INIT1 = 16'hf555;
    defparam add_1176_21.INJECT1_0 = "NO";
    defparam add_1176_21.INJECT1_1 = "NO";
    FD1P3IX intgOut2_i19 (.D(intgOut0_28__N_1433[19]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i19.GSR = "ENABLED";
    FD1P3IX intgOut2_i18 (.D(intgOut0_28__N_1433[18]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i18.GSR = "ENABLED";
    FD1P3IX intgOut2_i17 (.D(intgOut0_28__N_1433[17]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i17.GSR = "ENABLED";
    FD1P3IX intgOut2_i16 (.D(intgOut0_28__N_1433[16]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i16.GSR = "ENABLED";
    FD1P3IX intgOut2_i15 (.D(intgOut0_28__N_1433[15]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i15.GSR = "ENABLED";
    FD1P3IX intgOut2_i14 (.D(intgOut0_28__N_1433[14]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i14.GSR = "ENABLED";
    FD1P3IX intgOut2_i13 (.D(intgOut0_28__N_1433[13]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i13.GSR = "ENABLED";
    CCU2D sub_16_rep_4_add_2_7 (.A0(n4384), .B0(n11439), .C0(n5776), .D0(n16270), 
          .A1(n4383), .B1(n11439), .C1(n5778), .D1(n16270), .CIN(n18235), 
          .COUT(n18236), .S0(n4456), .S1(n4455));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_7.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_7.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_7.INJECT1_1 = "NO";
    FD1P3IX intgOut2_i12 (.D(intgOut0_28__N_1433[12]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i12.GSR = "ENABLED";
    FD1P3IX intgOut2_i11 (.D(intgOut0_28__N_1433[11]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i11.GSR = "ENABLED";
    FD1P3IX intgOut2_i10 (.D(intgOut0_28__N_1433[10]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i10.GSR = "ENABLED";
    CCU2D add_1176_19 (.A0(n5404), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5406), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18030), 
          .COUT(n18031), .S0(n2341[17]), .S1(n2341[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1176_19.INIT0 = 16'hf555;
    defparam add_1176_19.INIT1 = 16'hf555;
    defparam add_1176_19.INJECT1_0 = "NO";
    defparam add_1176_19.INJECT1_1 = "NO";
    FD1P3IX intgOut2_i9 (.D(intgOut0_28__N_1433[9]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i9.GSR = "ENABLED";
    FD1P3IX intgOut2_i8 (.D(intgOut0_28__N_1433[8]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i8.GSR = "ENABLED";
    FD1P3IX intgOut2_i7 (.D(intgOut0_28__N_1433[7]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i7.GSR = "ENABLED";
    FD1P3IX intgOut2_i6 (.D(intgOut0_28__N_1433[6]), .SP(clk_N_683_enable_331), 
            .CD(n14284), .CK(clk_N_683), .Q(intgOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i6.GSR = "ENABLED";
    FD1P3IX intgOut2_i5 (.D(addOut[5]), .SP(clk_N_683_enable_331), .CD(n14278), 
            .CK(clk_N_683), .Q(intgOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i5.GSR = "ENABLED";
    FD1P3IX intgOut2_i4 (.D(addOut[4]), .SP(clk_N_683_enable_331), .CD(n14278), 
            .CK(clk_N_683), .Q(intgOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i4.GSR = "ENABLED";
    FD1P3IX intgOut2_i3 (.D(addOut[3]), .SP(clk_N_683_enable_331), .CD(n14278), 
            .CK(clk_N_683), .Q(intgOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i3.GSR = "ENABLED";
    FD1P3IX intgOut2_i2 (.D(addOut[2]), .SP(clk_N_683_enable_331), .CD(n14278), 
            .CK(clk_N_683), .Q(intgOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i2.GSR = "ENABLED";
    FD1P3IX intgOut2_i1 (.D(addOut[1]), .SP(clk_N_683_enable_331), .CD(n14278), 
            .CK(clk_N_683), .Q(intgOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i1.GSR = "ENABLED";
    FD1P3IX intgOut1_i28 (.D(intgOut0_28__N_1433[28]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i28.GSR = "ENABLED";
    FD1P3IX intgOut1_i27 (.D(intgOut0_28__N_1433[27]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i27.GSR = "ENABLED";
    CCU2D add_15006_11 (.A0(speed_set_m1[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18312), .COUT(n18313));
    defparam add_15006_11.INIT0 = 16'hf555;
    defparam add_15006_11.INIT1 = 16'hf555;
    defparam add_15006_11.INJECT1_0 = "NO";
    defparam add_15006_11.INJECT1_1 = "NO";
    PFUMX mux_140_i29 (.BLUT(n551[28]), .ALUT(n671[28]), .C0(n20019), 
          .Z(addIn2_28__N_1375[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i26 (.D(intgOut0_28__N_1433[26]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i26.GSR = "ENABLED";
    FD1P3IX intgOut1_i25 (.D(intgOut0_28__N_1433[25]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i25.GSR = "ENABLED";
    PFUMX mux_137_i2 (.BLUT(n581[1]), .ALUT(intgOut3[1]), .C0(n21308), 
          .Z(n611[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_2_lut_rep_397 (.A(n22105), .B(ss[3]), .Z(n21378)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam i1_2_lut_rep_397.init = 16'hbbbb;
    FD1P3IX intgOut1_i24 (.D(intgOut0_28__N_1433[24]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i24.GSR = "ENABLED";
    FD1P3IX intgOut1_i23 (.D(intgOut0_28__N_1433[23]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i23.GSR = "ENABLED";
    PFUMX mux_137_i3 (.BLUT(n581[2]), .ALUT(intgOut3[2]), .C0(n21308), 
          .Z(n611[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i22 (.D(intgOut0_28__N_1433[22]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i22.GSR = "ENABLED";
    FD1P3IX intgOut1_i21 (.D(intgOut0_28__N_1433[21]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i21.GSR = "ENABLED";
    PFUMX mux_137_i4 (.BLUT(n581[3]), .ALUT(intgOut3[3]), .C0(n21308), 
          .Z(n611[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i20 (.D(intgOut0_28__N_1433[20]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i20.GSR = "ENABLED";
    FD1P3IX intgOut1_i19 (.D(intgOut0_28__N_1433[19]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i19.GSR = "ENABLED";
    PFUMX mux_137_i5 (.BLUT(n581[4]), .ALUT(intgOut3[4]), .C0(n21308), 
          .Z(n611[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i18 (.D(intgOut0_28__N_1433[18]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i18.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_361_3_lut (.A(n22105), .B(ss[3]), .C(ss[2]), .Z(n21342)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam i1_2_lut_rep_361_3_lut.init = 16'hfbfb;
    FD1P3IX intgOut1_i17 (.D(intgOut0_28__N_1433[17]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i17.GSR = "ENABLED";
    LUT4 mux_251_i6_3_lut_4_lut_3_lut (.A(n30_adj_2145), .B(n1349[15]), 
         .C(n2285[5]), .Z(n1531[5])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[25:42])
    defparam mux_251_i6_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FD1P3IX intgOut1_i16 (.D(intgOut0_28__N_1433[16]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i16.GSR = "ENABLED";
    FD1P3IX intgOut1_i15 (.D(intgOut0_28__N_1433[15]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i15.GSR = "ENABLED";
    FD1P3IX intgOut1_i14 (.D(intgOut0_28__N_1433[14]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i14.GSR = "ENABLED";
    FD1P3IX intgOut1_i13 (.D(intgOut0_28__N_1433[13]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i13.GSR = "ENABLED";
    FD1P3IX intgOut1_i12 (.D(intgOut0_28__N_1433[12]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i12.GSR = "ENABLED";
    LUT4 mux_251_i10_3_lut_4_lut_3_lut (.A(n30_adj_2145), .B(n1349[15]), 
         .C(n2285[9]), .Z(n1531[9])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[25:42])
    defparam mux_251_i10_3_lut_4_lut_3_lut.init = 16'hc4c4;
    PFUMX mux_137_i6 (.BLUT(n581[5]), .ALUT(intgOut3[5]), .C0(n21308), 
          .Z(n611[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i11 (.D(intgOut0_28__N_1433[11]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i11.GSR = "ENABLED";
    FD1P3IX intgOut1_i10 (.D(intgOut0_28__N_1433[10]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i10.GSR = "ENABLED";
    FD1P3IX intgOut1_i9 (.D(intgOut0_28__N_1433[9]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i9.GSR = "ENABLED";
    LUT4 mux_91_i4_3_lut_4_lut_4_lut (.A(n21308), .B(\speed_avg_m4[3] ), 
         .C(n4322), .D(n22082), .Z(n367[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i4_3_lut_4_lut_4_lut.init = 16'hcacf;
    FD1P3IX intgOut1_i8 (.D(intgOut0_28__N_1433[8]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i8.GSR = "ENABLED";
    LUT4 mux_251_i7_3_lut_4_lut_3_lut (.A(n30_adj_2145), .B(n1349[15]), 
         .C(n2285[6]), .Z(n1531[6])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[25:42])
    defparam mux_251_i7_3_lut_4_lut_3_lut.init = 16'hc4c4;
    PFUMX mux_137_i7 (.BLUT(n581[6]), .ALUT(intgOut3[6]), .C0(n21308), 
          .Z(n611[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i7 (.D(intgOut0_28__N_1433[7]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i7.GSR = "ENABLED";
    FD1P3IX intgOut1_i6 (.D(intgOut0_28__N_1433[6]), .SP(clk_N_683_enable_390), 
            .CD(n14256), .CK(clk_N_683), .Q(intgOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i6.GSR = "ENABLED";
    FD1P3IX intgOut1_i5 (.D(addOut[5]), .SP(clk_N_683_enable_390), .CD(n14250), 
            .CK(clk_N_683), .Q(intgOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i5.GSR = "ENABLED";
    FD1P3IX intgOut1_i4 (.D(addOut[4]), .SP(clk_N_683_enable_390), .CD(n14250), 
            .CK(clk_N_683), .Q(intgOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i4.GSR = "ENABLED";
    PFUMX mux_137_i8 (.BLUT(n581[7]), .ALUT(intgOut3[7]), .C0(n21308), 
          .Z(n611[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i9 (.BLUT(n581[8]), .ALUT(intgOut3[8]), .C0(n21308), 
          .Z(n611[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut1_i3 (.D(addOut[3]), .SP(clk_N_683_enable_390), .CD(n14250), 
            .CK(clk_N_683), .Q(intgOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i3.GSR = "ENABLED";
    FD1P3IX intgOut1_i2 (.D(addOut[2]), .SP(clk_N_683_enable_390), .CD(n14250), 
            .CK(clk_N_683), .Q(intgOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i2.GSR = "ENABLED";
    FD1P3IX intgOut1_i1 (.D(addOut[1]), .SP(clk_N_683_enable_390), .CD(n14250), 
            .CK(clk_N_683), .Q(intgOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i1.GSR = "ENABLED";
    PFUMX mux_137_i10 (.BLUT(n581[9]), .ALUT(intgOut3[9]), .C0(n21308), 
          .Z(n611[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i28 (.D(intgOut0_28__N_1433[28]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i28.GSR = "ENABLED";
    PFUMX mux_137_i11 (.BLUT(n581[10]), .ALUT(intgOut3[10]), .C0(n21308), 
          .Z(n611[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 ss_4__I_0_355_i9_2_lut_3_lut_4_lut (.A(n22105), .B(ss[3]), .C(n21379), 
         .D(n22099), .Z(n9_adj_2137)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam ss_4__I_0_355_i9_2_lut_3_lut_4_lut.init = 16'hfffb;
    FD1P3IX intgOut0_i27 (.D(intgOut0_28__N_1433[27]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i27.GSR = "ENABLED";
    FD1P3IX intgOut0_i26 (.D(intgOut0_28__N_1433[26]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i26.GSR = "ENABLED";
    FD1P3IX intgOut0_i25 (.D(intgOut0_28__N_1433[25]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i25.GSR = "ENABLED";
    LUT4 mux_251_i8_3_lut_4_lut_3_lut (.A(n30_adj_2145), .B(n1349[15]), 
         .C(n2285[7]), .Z(n1531[7])) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[25:42])
    defparam mux_251_i8_3_lut_4_lut_3_lut.init = 16'hc4c4;
    FD1P3IX intgOut0_i24 (.D(intgOut0_28__N_1433[24]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i24.GSR = "ENABLED";
    FD1P3IX intgOut0_i23 (.D(intgOut0_28__N_1433[23]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i23.GSR = "ENABLED";
    FD1P3IX intgOut0_i22 (.D(intgOut0_28__N_1433[22]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i22.GSR = "ENABLED";
    FD1P3IX intgOut0_i21 (.D(intgOut0_28__N_1433[21]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i21.GSR = "ENABLED";
    PFUMX mux_137_i12 (.BLUT(n581[11]), .ALUT(intgOut3[11]), .C0(n21308), 
          .Z(n611[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i20 (.D(intgOut0_28__N_1433[20]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i20.GSR = "ENABLED";
    FD1P3IX intgOut0_i19 (.D(intgOut0_28__N_1433[19]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i19.GSR = "ENABLED";
    FD1P3IX intgOut0_i18 (.D(intgOut0_28__N_1433[18]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i18.GSR = "ENABLED";
    FD1P3IX intgOut0_i17 (.D(intgOut0_28__N_1433[17]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i17.GSR = "ENABLED";
    LUT4 equal_112_i9_2_lut_3_lut_4_lut (.A(n22105), .B(ss[3]), .C(n21379), 
         .D(ss[2]), .Z(n9_adj_2138)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam equal_112_i9_2_lut_3_lut_4_lut.init = 16'hfbff;
    FD1P3IX intgOut0_i16 (.D(intgOut0_28__N_1433[16]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i16.GSR = "ENABLED";
    PFUMX mux_137_i13 (.BLUT(n581[12]), .ALUT(intgOut3[12]), .C0(n21308), 
          .Z(n611[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i15 (.D(intgOut0_28__N_1433[15]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i15.GSR = "ENABLED";
    FD1P3IX intgOut0_i14 (.D(intgOut0_28__N_1433[14]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i14.GSR = "ENABLED";
    LUT4 i13380_2_lut (.A(addOut[18]), .B(n22105), .Z(backOut3_28__N_1678[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13380_2_lut.init = 16'h2222;
    FD1P3IX intgOut0_i13 (.D(intgOut0_28__N_1433[13]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i13.GSR = "ENABLED";
    LUT4 ss_4__I_0_355_i6_2_lut_rep_398 (.A(ss[0]), .B(ss[1]), .Z(n21379)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(167[9:16])
    defparam ss_4__I_0_355_i6_2_lut_rep_398.init = 16'heeee;
    PFUMX mux_137_i14 (.BLUT(n581[13]), .ALUT(intgOut3[13]), .C0(n21308), 
          .Z(n611[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i12 (.D(intgOut0_28__N_1433[12]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i12.GSR = "ENABLED";
    FD1P3IX intgOut0_i11 (.D(intgOut0_28__N_1433[11]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i11.GSR = "ENABLED";
    CCU2D add_15006_9 (.A0(speed_set_m1[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18311), .COUT(n18312));
    defparam add_15006_9.INIT0 = 16'hf555;
    defparam add_15006_9.INIT1 = 16'hf555;
    defparam add_15006_9.INJECT1_0 = "NO";
    defparam add_15006_9.INJECT1_1 = "NO";
    FD1P3IX intgOut0_i10 (.D(intgOut0_28__N_1433[10]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i10.GSR = "ENABLED";
    LUT4 i2_4_lut_then_3_lut (.A(ss[0]), .B(n21342), .C(n21325), .Z(n22094)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i2_4_lut_then_3_lut.init = 16'he0e0;
    FD1P3IX intgOut0_i9 (.D(intgOut0_28__N_1433[9]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i9.GSR = "ENABLED";
    FD1P3IX intgOut0_i8 (.D(intgOut0_28__N_1433[8]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i8.GSR = "ENABLED";
    PFUMX mux_137_i15 (.BLUT(n581[14]), .ALUT(intgOut3[14]), .C0(n21308), 
          .Z(n611[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i7 (.D(intgOut0_28__N_1433[7]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i7.GSR = "ENABLED";
    FD1P3IX intgOut0_i6 (.D(intgOut0_28__N_1433[6]), .SP(clk_N_683_enable_387), 
            .CD(n14228), .CK(clk_N_683), .Q(intgOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i6.GSR = "ENABLED";
    FD1P3IX intgOut0_i5 (.D(addOut[5]), .SP(clk_N_683_enable_387), .CD(n14222), 
            .CK(clk_N_683), .Q(intgOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i5.GSR = "ENABLED";
    PFUMX mux_137_i16 (.BLUT(n581[15]), .ALUT(intgOut3[15]), .C0(n21308), 
          .Z(n611[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    FD1P3IX intgOut0_i4 (.D(addOut[4]), .SP(clk_N_683_enable_387), .CD(n14222), 
            .CK(clk_N_683), .Q(intgOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i4.GSR = "ENABLED";
    FD1P3IX intgOut0_i3 (.D(addOut[3]), .SP(clk_N_683_enable_387), .CD(n14222), 
            .CK(clk_N_683), .Q(intgOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i3.GSR = "ENABLED";
    FD1P3IX intgOut0_i2 (.D(addOut[2]), .SP(clk_N_683_enable_387), .CD(n14222), 
            .CK(clk_N_683), .Q(intgOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i2.GSR = "ENABLED";
    FD1P3IX intgOut0_i1 (.D(addOut[1]), .SP(clk_N_683_enable_387), .CD(n14222), 
            .CK(clk_N_683), .Q(intgOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i1.GSR = "ENABLED";
    PFUMX mux_137_i17 (.BLUT(n581[16]), .ALUT(intgOut3[16]), .C0(n21308), 
          .Z(n611[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D sub_16_rep_4_add_2_5 (.A0(n4386), .B0(n11439), .C0(n5772), .D0(n16270), 
          .A1(n4385), .B1(n11439), .C1(n5774), .D1(n16270), .CIN(n18234), 
          .COUT(n18235), .S0(n4458), .S1(n4457));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_5.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_5.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_5.INJECT1_1 = "NO";
    LUT4 ss_4__I_0_357_i9_2_lut_rep_344_3_lut_4_lut (.A(n22105), .B(ss[3]), 
         .C(n22083), .D(ss[2]), .Z(n21325)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam ss_4__I_0_357_i9_2_lut_rep_344_3_lut_4_lut.init = 16'hffef;
    CCU2D add_15006_7 (.A0(speed_set_m1[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18310), .COUT(n18311));
    defparam add_15006_7.INIT0 = 16'hf555;
    defparam add_15006_7.INIT1 = 16'hf555;
    defparam add_15006_7.INJECT1_0 = "NO";
    defparam add_15006_7.INJECT1_1 = "NO";
    CCU2D add_1173_11 (.A0(n1349[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18149), 
          .S0(n2285[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1173_11.INIT0 = 16'hf555;
    defparam add_1173_11.INIT1 = 16'h0000;
    defparam add_1173_11.INJECT1_0 = "NO";
    defparam add_1173_11.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_3 (.A0(n4388), .B0(n11439), .C0(n5768), .D0(n16270), 
          .A1(n4387), .B1(n11439), .C1(n5770), .D1(n16270), .CIN(n18233), 
          .COUT(n18234), .S0(n4460), .S1(n4459));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_3.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_3.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n4389), .B1(n11439), .C1(n5481), .D1(n16270), 
          .COUT(n18233), .S1(n4461));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_1.INIT0 = 16'h0000;
    defparam sub_16_rep_4_add_2_1.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_1.INJECT1_1 = "NO";
    CCU2D add_1173_9 (.A0(n1349[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1349[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18148), 
          .COUT(n18149), .S0(n2285[7]), .S1(n2285[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1173_9.INIT0 = 16'hf555;
    defparam add_1173_9.INIT1 = 16'hf555;
    defparam add_1173_9.INJECT1_0 = "NO";
    defparam add_1173_9.INJECT1_1 = "NO";
    CCU2D add_15006_5 (.A0(speed_set_m1[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18309), .COUT(n18310));
    defparam add_15006_5.INIT0 = 16'hf555;
    defparam add_15006_5.INIT1 = 16'hf555;
    defparam add_15006_5.INJECT1_0 = "NO";
    defparam add_15006_5.INJECT1_1 = "NO";
    CCU2D add_15006_3 (.A0(speed_set_m1[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18308), .COUT(n18309));
    defparam add_15006_3.INIT0 = 16'hf555;
    defparam add_15006_3.INIT1 = 16'hf555;
    defparam add_15006_3.INJECT1_0 = "NO";
    defparam add_15006_3.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_29 (.A0(multOut[27]), .B0(n16396), .C0(addOut[27]), 
          .D0(addIn2_28__N_1246[27]), .A1(multOut[28]), .B1(n16396), .C1(addOut[28]), 
          .D1(addIn2_28__N_1246[28]), .CIN(n18231), .S0(n121[27]), .S1(n121[28]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_29.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_29.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_29.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_29.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_360_3_lut (.A(n22105), .B(ss[3]), .C(n22099), .Z(n21341)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_360_3_lut.init = 16'hfefe;
    CCU2D add_15006_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[0]), .B1(speed_set_m1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18308));
    defparam add_15006_1.INIT0 = 16'hF000;
    defparam add_15006_1.INIT1 = 16'ha666;
    defparam add_15006_1.INJECT1_0 = "NO";
    defparam add_15006_1.INJECT1_1 = "NO";
    CCU2D add_1173_7 (.A0(n1349[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1349[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18147), 
          .COUT(n18148), .S0(n2285[5]), .S1(n2285[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1173_7.INIT0 = 16'hf555;
    defparam add_1173_7.INIT1 = 16'hf555;
    defparam add_1173_7.INJECT1_0 = "NO";
    defparam add_1173_7.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_27 (.A0(multOut[25]), .B0(n16396), .C0(addOut[25]), 
          .D0(addIn2_28__N_1246[25]), .A1(multOut[26]), .B1(n16396), .C1(addOut[26]), 
          .D1(addIn2_28__N_1246[26]), .CIN(n18230), .COUT(n18231), .S0(n121[25]), 
          .S1(n121[26]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_27.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_27.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_27.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_27.INJECT1_1 = "NO";
    PFUMX mux_137_i18 (.BLUT(n581[17]), .ALUT(intgOut3[17]), .C0(n21308), 
          .Z(n611[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i19 (.BLUT(n581[18]), .ALUT(intgOut3[18]), .C0(n21308), 
          .Z(n611[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i20 (.BLUT(n581[19]), .ALUT(intgOut3[19]), .C0(n21308), 
          .Z(n611[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i21 (.BLUT(n581[20]), .ALUT(intgOut3[20]), .C0(n21308), 
          .Z(n611[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i22 (.BLUT(n581[21]), .ALUT(intgOut3[21]), .C0(n21308), 
          .Z(n611[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_2_lut_rep_363_3_lut (.A(n22105), .B(ss[3]), .C(n22099), .Z(n21344)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_363_3_lut.init = 16'hefef;
    PFUMX mux_137_i23 (.BLUT(n581[22]), .ALUT(intgOut3[22]), .C0(n21308), 
          .Z(n611[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    PFUMX mux_137_i24 (.BLUT(n581[23]), .ALUT(intgOut3[23]), .C0(n21308), 
          .Z(n611[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i7911_2_lut_3_lut (.A(ss[0]), .B(ss[1]), .C(ss[2]), .Z(n14)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i7911_2_lut_3_lut.init = 16'h7878;
    PFUMX mux_137_i25 (.BLUT(n581[24]), .ALUT(intgOut3[24]), .C0(n21308), 
          .Z(n611[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i1_2_lut_rep_365_3_lut_4_lut (.A(n22105), .B(ss[3]), .C(ss[1]), 
         .D(ss[0]), .Z(n21346)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_rep_365_3_lut_4_lut.init = 16'h0110;
    PFUMX mux_137_i26 (.BLUT(n581[25]), .ALUT(intgOut3[25]), .C0(n21308), 
          .Z(n611[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_14994_17 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18434), .S1(n3744));
    defparam add_14994_17.INIT0 = 16'h5555;
    defparam add_14994_17.INIT1 = 16'h0000;
    defparam add_14994_17.INJECT1_0 = "NO";
    defparam add_14994_17.INJECT1_1 = "NO";
    LUT4 i16252_2_lut_rep_401 (.A(ss[2]), .B(ss[3]), .Z(n21382)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16252_2_lut_rep_401.init = 16'h8888;
    CCU2D add_14994_15 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18433), .COUT(n18434));
    defparam add_14994_15.INIT0 = 16'hf555;
    defparam add_14994_15.INIT1 = 16'hf555;
    defparam add_14994_15.INJECT1_0 = "NO";
    defparam add_14994_15.INJECT1_1 = "NO";
    CCU2D add_14994_13 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18432), .COUT(n18433));
    defparam add_14994_13.INIT0 = 16'hf555;
    defparam add_14994_13.INIT1 = 16'hf555;
    defparam add_14994_13.INJECT1_0 = "NO";
    defparam add_14994_13.INJECT1_1 = "NO";
    CCU2D add_14994_11 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18431), .COUT(n18432));
    defparam add_14994_11.INIT0 = 16'hf555;
    defparam add_14994_11.INIT1 = 16'hf555;
    defparam add_14994_11.INJECT1_0 = "NO";
    defparam add_14994_11.INJECT1_1 = "NO";
    CCU2D add_14994_9 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18430), .COUT(n18431));
    defparam add_14994_9.INIT0 = 16'hf555;
    defparam add_14994_9.INIT1 = 16'h0aaa;
    defparam add_14994_9.INJECT1_0 = "NO";
    defparam add_14994_9.INJECT1_1 = "NO";
    CCU2D add_14994_7 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18429), .COUT(n18430));
    defparam add_14994_7.INIT0 = 16'h0aaa;
    defparam add_14994_7.INIT1 = 16'hf555;
    defparam add_14994_7.INJECT1_0 = "NO";
    defparam add_14994_7.INJECT1_1 = "NO";
    LUT4 ss_4__I_0_360_i9_2_lut_rep_345_3_lut_4_lut (.A(n22105), .B(ss[3]), 
         .C(n22083), .D(ss[2]), .Z(n21326)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam ss_4__I_0_360_i9_2_lut_rep_345_3_lut_4_lut.init = 16'hefff;
    LUT4 ss_1__bdd_3_lut_4_lut (.A(ss[2]), .B(ss[3]), .C(ss[0]), .D(ss[1]), 
         .Z(n21243)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam ss_1__bdd_3_lut_4_lut.init = 16'h0800;
    CCU2D add_14994_5 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18428), .COUT(n18429));
    defparam add_14994_5.INIT0 = 16'h0aaa;
    defparam add_14994_5.INIT1 = 16'h0aaa;
    defparam add_14994_5.INJECT1_0 = "NO";
    defparam add_14994_5.INJECT1_1 = "NO";
    CCU2D add_14994_3 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18427), .COUT(n18428));
    defparam add_14994_3.INIT0 = 16'hf555;
    defparam add_14994_3.INIT1 = 16'hf555;
    defparam add_14994_3.INJECT1_0 = "NO";
    defparam add_14994_3.INJECT1_1 = "NO";
    CCU2D add_14994_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[4]), .B1(speed_set_m4[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18427));
    defparam add_14994_1.INIT0 = 16'hF000;
    defparam add_14994_1.INIT1 = 16'ha666;
    defparam add_14994_1.INJECT1_0 = "NO";
    defparam add_14994_1.INJECT1_1 = "NO";
    CCU2D add_14995_29 (.A0(addOut[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18426), 
          .S1(n3832));
    defparam add_14995_29.INIT0 = 16'h5aaa;
    defparam add_14995_29.INIT1 = 16'h0000;
    defparam add_14995_29.INJECT1_0 = "NO";
    defparam add_14995_29.INJECT1_1 = "NO";
    CCU2D add_14995_27 (.A0(addOut[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18425), .COUT(n18426));
    defparam add_14995_27.INIT0 = 16'h0aaa;
    defparam add_14995_27.INIT1 = 16'h0aaa;
    defparam add_14995_27.INJECT1_0 = "NO";
    defparam add_14995_27.INJECT1_1 = "NO";
    CCU2D add_14995_25 (.A0(addOut[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18424), .COUT(n18425));
    defparam add_14995_25.INIT0 = 16'h0aaa;
    defparam add_14995_25.INIT1 = 16'h0aaa;
    defparam add_14995_25.INJECT1_0 = "NO";
    defparam add_14995_25.INJECT1_1 = "NO";
    CCU2D add_14995_23 (.A0(addOut[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18423), .COUT(n18424));
    defparam add_14995_23.INIT0 = 16'h0aaa;
    defparam add_14995_23.INIT1 = 16'h0aaa;
    defparam add_14995_23.INJECT1_0 = "NO";
    defparam add_14995_23.INJECT1_1 = "NO";
    CCU2D add_14995_21 (.A0(addOut[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18422), .COUT(n18423));
    defparam add_14995_21.INIT0 = 16'h0aaa;
    defparam add_14995_21.INIT1 = 16'h0aaa;
    defparam add_14995_21.INJECT1_0 = "NO";
    defparam add_14995_21.INJECT1_1 = "NO";
    CCU2D add_14995_19 (.A0(addOut[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18421), .COUT(n18422));
    defparam add_14995_19.INIT0 = 16'hf555;
    defparam add_14995_19.INIT1 = 16'hf555;
    defparam add_14995_19.INJECT1_0 = "NO";
    defparam add_14995_19.INJECT1_1 = "NO";
    CCU2D add_14995_17 (.A0(addOut[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18420), .COUT(n18421));
    defparam add_14995_17.INIT0 = 16'hf555;
    defparam add_14995_17.INIT1 = 16'hf555;
    defparam add_14995_17.INJECT1_0 = "NO";
    defparam add_14995_17.INJECT1_1 = "NO";
    CCU2D add_14995_15 (.A0(addOut[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18419), .COUT(n18420));
    defparam add_14995_15.INIT0 = 16'hf555;
    defparam add_14995_15.INIT1 = 16'h0aaa;
    defparam add_14995_15.INJECT1_0 = "NO";
    defparam add_14995_15.INJECT1_1 = "NO";
    CCU2D add_14995_13 (.A0(addOut[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18418), .COUT(n18419));
    defparam add_14995_13.INIT0 = 16'h0aaa;
    defparam add_14995_13.INIT1 = 16'h0aaa;
    defparam add_14995_13.INJECT1_0 = "NO";
    defparam add_14995_13.INJECT1_1 = "NO";
    CCU2D add_14995_11 (.A0(addOut[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18417), .COUT(n18418));
    defparam add_14995_11.INIT0 = 16'h0aaa;
    defparam add_14995_11.INIT1 = 16'h0aaa;
    defparam add_14995_11.INJECT1_0 = "NO";
    defparam add_14995_11.INJECT1_1 = "NO";
    CCU2D add_14995_9 (.A0(addOut[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18416), .COUT(n18417));
    defparam add_14995_9.INIT0 = 16'h0aaa;
    defparam add_14995_9.INIT1 = 16'hf555;
    defparam add_14995_9.INJECT1_0 = "NO";
    defparam add_14995_9.INJECT1_1 = "NO";
    CCU2D add_14995_7 (.A0(addOut[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18415), .COUT(n18416));
    defparam add_14995_7.INIT0 = 16'h0aaa;
    defparam add_14995_7.INIT1 = 16'h0aaa;
    defparam add_14995_7.INJECT1_0 = "NO";
    defparam add_14995_7.INJECT1_1 = "NO";
    LUT4 i13373_2_lut (.A(addOut[17]), .B(n22105), .Z(backOut3_28__N_1678[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13373_2_lut.init = 16'h2222;
    CCU2D add_14995_5 (.A0(addOut[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18414), .COUT(n18415));
    defparam add_14995_5.INIT0 = 16'hf555;
    defparam add_14995_5.INIT1 = 16'hf555;
    defparam add_14995_5.INJECT1_0 = "NO";
    defparam add_14995_5.INJECT1_1 = "NO";
    PFUMX mux_137_i27 (.BLUT(n581[26]), .ALUT(intgOut3[26]), .C0(n21308), 
          .Z(n611[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_14995_3 (.A0(addOut[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18413), .COUT(n18414));
    defparam add_14995_3.INIT0 = 16'hf555;
    defparam add_14995_3.INIT1 = 16'hf555;
    defparam add_14995_3.INJECT1_0 = "NO";
    defparam add_14995_3.INJECT1_1 = "NO";
    CCU2D add_14995_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[0]), .B1(addOut[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18413));
    defparam add_14995_1.INIT0 = 16'hF000;
    defparam add_14995_1.INIT1 = 16'ha666;
    defparam add_14995_1.INJECT1_0 = "NO";
    defparam add_14995_1.INJECT1_1 = "NO";
    CCU2D add_14996_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18412), 
          .S0(n1061));
    defparam add_14996_cout.INIT0 = 16'h0000;
    defparam add_14996_cout.INIT1 = 16'h0000;
    defparam add_14996_cout.INJECT1_0 = "NO";
    defparam add_14996_cout.INJECT1_1 = "NO";
    CCU2D add_14996_22 (.A0(addOut[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18411), .COUT(n18412));
    defparam add_14996_22.INIT0 = 16'h5555;
    defparam add_14996_22.INIT1 = 16'hf555;
    defparam add_14996_22.INJECT1_0 = "NO";
    defparam add_14996_22.INJECT1_1 = "NO";
    CCU2D add_14996_20 (.A0(addOut[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18410), .COUT(n18411));
    defparam add_14996_20.INIT0 = 16'h5555;
    defparam add_14996_20.INIT1 = 16'h5555;
    defparam add_14996_20.INJECT1_0 = "NO";
    defparam add_14996_20.INJECT1_1 = "NO";
    CCU2D add_14996_18 (.A0(addOut[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18409), .COUT(n18410));
    defparam add_14996_18.INIT0 = 16'h5555;
    defparam add_14996_18.INIT1 = 16'h5555;
    defparam add_14996_18.INJECT1_0 = "NO";
    defparam add_14996_18.INJECT1_1 = "NO";
    CCU2D add_14996_16 (.A0(addOut[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18408), .COUT(n18409));
    defparam add_14996_16.INIT0 = 16'h5555;
    defparam add_14996_16.INIT1 = 16'h5555;
    defparam add_14996_16.INJECT1_0 = "NO";
    defparam add_14996_16.INJECT1_1 = "NO";
    CCU2D add_14996_14 (.A0(addOut[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18407), .COUT(n18408));
    defparam add_14996_14.INIT0 = 16'h5aaa;
    defparam add_14996_14.INIT1 = 16'h5555;
    defparam add_14996_14.INJECT1_0 = "NO";
    defparam add_14996_14.INJECT1_1 = "NO";
    LUT4 i13367_2_lut (.A(addOut[15]), .B(n22105), .Z(backOut3_28__N_1678[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13367_2_lut.init = 16'h2222;
    CCU2D add_14996_12 (.A0(addOut[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18406), .COUT(n18407));
    defparam add_14996_12.INIT0 = 16'h5aaa;
    defparam add_14996_12.INIT1 = 16'h5aaa;
    defparam add_14996_12.INJECT1_0 = "NO";
    defparam add_14996_12.INJECT1_1 = "NO";
    CCU2D add_14996_10 (.A0(addOut[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18405), .COUT(n18406));
    defparam add_14996_10.INIT0 = 16'h5555;
    defparam add_14996_10.INIT1 = 16'h5aaa;
    defparam add_14996_10.INJECT1_0 = "NO";
    defparam add_14996_10.INJECT1_1 = "NO";
    CCU2D add_14996_8 (.A0(addOut[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18404), .COUT(n18405));
    defparam add_14996_8.INIT0 = 16'h5555;
    defparam add_14996_8.INIT1 = 16'h5aaa;
    defparam add_14996_8.INJECT1_0 = "NO";
    defparam add_14996_8.INJECT1_1 = "NO";
    CCU2D add_14996_6 (.A0(addOut[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18403), .COUT(n18404));
    defparam add_14996_6.INIT0 = 16'h5555;
    defparam add_14996_6.INIT1 = 16'h5555;
    defparam add_14996_6.INJECT1_0 = "NO";
    defparam add_14996_6.INJECT1_1 = "NO";
    CCU2D add_14996_4 (.A0(addOut[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18402), .COUT(n18403));
    defparam add_14996_4.INIT0 = 16'h5aaa;
    defparam add_14996_4.INIT1 = 16'h5555;
    defparam add_14996_4.INJECT1_0 = "NO";
    defparam add_14996_4.INJECT1_1 = "NO";
    CCU2D add_14996_2 (.A0(addOut[7]), .B0(addOut[6]), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18402));
    defparam add_14996_2.INIT0 = 16'h1000;
    defparam add_14996_2.INIT1 = 16'h5555;
    defparam add_14996_2.INJECT1_0 = "NO";
    defparam add_14996_2.INJECT1_1 = "NO";
    CCU2D add_14997_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18401), 
          .S0(n3768));
    defparam add_14997_cout.INIT0 = 16'h0000;
    defparam add_14997_cout.INIT1 = 16'h0000;
    defparam add_14997_cout.INJECT1_0 = "NO";
    defparam add_14997_cout.INJECT1_1 = "NO";
    CCU2D add_14997_20 (.A0(speed_set_m4[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18400), .COUT(n18401));
    defparam add_14997_20.INIT0 = 16'h5aaa;
    defparam add_14997_20.INIT1 = 16'h0aaa;
    defparam add_14997_20.INJECT1_0 = "NO";
    defparam add_14997_20.INJECT1_1 = "NO";
    LUT4 mux_189_i20_3_lut_3_lut (.A(n1061), .B(n3832), .C(addOut[19]), 
         .Z(intgOut0_28__N_1433[19])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i20_3_lut_3_lut.init = 16'hbaba;
    CCU2D add_14997_18 (.A0(speed_set_m4[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18399), .COUT(n18400));
    defparam add_14997_18.INIT0 = 16'h5aaa;
    defparam add_14997_18.INIT1 = 16'h5aaa;
    defparam add_14997_18.INJECT1_0 = "NO";
    defparam add_14997_18.INJECT1_1 = "NO";
    CCU2D add_14997_16 (.A0(speed_set_m4[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18398), .COUT(n18399));
    defparam add_14997_16.INIT0 = 16'h5aaa;
    defparam add_14997_16.INIT1 = 16'h5aaa;
    defparam add_14997_16.INJECT1_0 = "NO";
    defparam add_14997_16.INJECT1_1 = "NO";
    CCU2D add_14997_14 (.A0(speed_set_m4[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18397), .COUT(n18398));
    defparam add_14997_14.INIT0 = 16'h5555;
    defparam add_14997_14.INIT1 = 16'h5aaa;
    defparam add_14997_14.INJECT1_0 = "NO";
    defparam add_14997_14.INJECT1_1 = "NO";
    CCU2D add_14997_12 (.A0(speed_set_m4[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18396), .COUT(n18397));
    defparam add_14997_12.INIT0 = 16'h5aaa;
    defparam add_14997_12.INIT1 = 16'h5aaa;
    defparam add_14997_12.INJECT1_0 = "NO";
    defparam add_14997_12.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_25 (.A0(multOut[23]), .B0(n16396), .C0(addOut[23]), 
          .D0(addIn2_28__N_1246[23]), .A1(multOut[24]), .B1(n16396), .C1(addOut[24]), 
          .D1(addIn2_28__N_1246[24]), .CIN(n18229), .COUT(n18230), .S0(n121[23]), 
          .S1(n121[24]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_25.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_25.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_25.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_25.INJECT1_1 = "NO";
    CCU2D add_14997_10 (.A0(speed_set_m4[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18395), .COUT(n18396));
    defparam add_14997_10.INIT0 = 16'h5555;
    defparam add_14997_10.INIT1 = 16'h5555;
    defparam add_14997_10.INJECT1_0 = "NO";
    defparam add_14997_10.INJECT1_1 = "NO";
    CCU2D add_1173_5 (.A0(n1349[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1349[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18146), 
          .COUT(n18147), .S0(n2285[3]), .S1(n2285[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1173_5.INIT0 = 16'hf555;
    defparam add_1173_5.INIT1 = 16'hf555;
    defparam add_1173_5.INJECT1_0 = "NO";
    defparam add_1173_5.INJECT1_1 = "NO";
    CCU2D add_1173_3 (.A0(n1349[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1349[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18145), 
          .COUT(n18146), .S0(n2285[1]), .S1(n2285[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1173_3.INIT0 = 16'hf555;
    defparam add_1173_3.INIT1 = 16'hf555;
    defparam add_1173_3.INJECT1_0 = "NO";
    defparam add_1173_3.INJECT1_1 = "NO";
    CCU2D add_14997_8 (.A0(speed_set_m4[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18394), .COUT(n18395));
    defparam add_14997_8.INIT0 = 16'h5aaa;
    defparam add_14997_8.INIT1 = 16'h5555;
    defparam add_14997_8.INJECT1_0 = "NO";
    defparam add_14997_8.INJECT1_1 = "NO";
    CCU2D add_1173_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1349[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18145), 
          .S1(n2285[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1173_1.INIT0 = 16'hF000;
    defparam add_1173_1.INIT1 = 16'h0aaa;
    defparam add_1173_1.INJECT1_0 = "NO";
    defparam add_1173_1.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_23 (.A0(multOut[21]), .B0(n16396), .C0(addOut[21]), 
          .D0(addIn2_28__N_1246[21]), .A1(multOut[22]), .B1(n16396), .C1(addOut[22]), 
          .D1(addIn2_28__N_1246[22]), .CIN(n18228), .COUT(n18229), .S0(n121[21]), 
          .S1(n121[22]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_23.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_23.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_23.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_23.INJECT1_1 = "NO";
    CCU2D add_14997_6 (.A0(speed_set_m4[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18393), .COUT(n18394));
    defparam add_14997_6.INIT0 = 16'h5aaa;
    defparam add_14997_6.INIT1 = 16'h5aaa;
    defparam add_14997_6.INJECT1_0 = "NO";
    defparam add_14997_6.INJECT1_1 = "NO";
    LUT4 i11538_3_lut_4_lut (.A(n1061), .B(n3832), .C(n21312), .D(clk_N_683_enable_303), 
         .Z(n14307)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i11538_3_lut_4_lut.init = 16'hfe00;
    CCU2D addOut_2081_add_4_21 (.A0(multOut[19]), .B0(n16396), .C0(addOut[19]), 
          .D0(addIn2_28__N_1246[19]), .A1(multOut[20]), .B1(n16396), .C1(addOut[20]), 
          .D1(addIn2_28__N_1246[20]), .CIN(n18227), .COUT(n18228), .S0(n121[19]), 
          .S1(n121[20]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_21.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_21.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_21.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_21.INJECT1_1 = "NO";
    CCU2D add_14997_4 (.A0(speed_set_m4[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18392), .COUT(n18393));
    defparam add_14997_4.INIT0 = 16'h5555;
    defparam add_14997_4.INIT1 = 16'h5aaa;
    defparam add_14997_4.INJECT1_0 = "NO";
    defparam add_14997_4.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_19 (.A0(multOut[17]), .B0(n16396), .C0(addOut[17]), 
          .D0(addIn2_28__N_1246[17]), .A1(multOut[18]), .B1(n16396), .C1(addOut[18]), 
          .D1(addIn2_28__N_1246[18]), .CIN(n18226), .COUT(n18227), .S0(n121[17]), 
          .S1(n121[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_19.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_19.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_19.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_19.INJECT1_1 = "NO";
    CCU2D add_1172_11 (.A0(n1328[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18144), 
          .S0(n2273[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1172_11.INIT0 = 16'hf555;
    defparam add_1172_11.INIT1 = 16'h0000;
    defparam add_1172_11.INJECT1_0 = "NO";
    defparam add_1172_11.INJECT1_1 = "NO";
    CCU2D add_14997_2 (.A0(speed_set_m4[1]), .B0(speed_set_m4[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18392));
    defparam add_14997_2.INIT0 = 16'h1000;
    defparam add_14997_2.INIT1 = 16'h5555;
    defparam add_14997_2.INJECT1_0 = "NO";
    defparam add_14997_2.INJECT1_1 = "NO";
    PFUMX mux_137_i28 (.BLUT(n581[27]), .ALUT(intgOut3[27]), .C0(n21308), 
          .Z(n611[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 i13364_2_lut (.A(addOut[14]), .B(n22105), .Z(backOut3_28__N_1678[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13364_2_lut.init = 16'h2222;
    LUT4 i13363_2_lut (.A(addOut[13]), .B(n22105), .Z(backOut3_28__N_1678[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13363_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(ss[2]), .B(n22105), .C(ss[3]), 
         .D(ss[0]), .Z(n16396)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(166[9:16])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hffed;
    LUT4 i17093_3_lut_3_lut_4_lut_4_lut_4_lut (.A(ss[0]), .B(n21344), .C(n21325), 
         .Z(n20019)) /* synthesis lut_function=(!(A (B (C))+!A (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(170[9:16])
    defparam i17093_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h2f2f;
    LUT4 i13362_2_lut (.A(addOut[12]), .B(n22105), .Z(backOut3_28__N_1678[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13362_2_lut.init = 16'h2222;
    LUT4 mux_1241_i6_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[5]), 
         .D(speed_set_m4[5]), .Z(n2581[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 i16644_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut (.A(ss[0]), .B(n21342), 
         .C(n9_adj_2138), .Z(n20022)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam i16644_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hd0d0;
    LUT4 ss_3__bdd_4_lut_17485 (.A(ss[3]), .B(n22105), .C(ss[1]), .D(ss[2]), 
         .Z(multIn2[4])) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam ss_3__bdd_4_lut_17485.init = 16'h0220;
    LUT4 i13361_2_lut (.A(addOut[11]), .B(n22105), .Z(backOut3_28__N_1678[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13361_2_lut.init = 16'h2222;
    CCU2D add_1172_9 (.A0(n1328[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1328[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18143), 
          .COUT(n18144), .S0(n2273[7]), .S1(n2273[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1172_9.INIT0 = 16'hf555;
    defparam add_1172_9.INIT1 = 16'hf555;
    defparam add_1172_9.INJECT1_0 = "NO";
    defparam add_1172_9.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_17 (.A0(multOut[15]), .B0(n16396), .C0(addOut[15]), 
          .D0(addIn2_28__N_1246[15]), .A1(multOut[16]), .B1(n16396), .C1(addOut[16]), 
          .D1(addIn2_28__N_1246[16]), .CIN(n18225), .COUT(n18226), .S0(n121[15]), 
          .S1(n121[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_17.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_17.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_17.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_17.INJECT1_1 = "NO";
    FD1P3IX dutyout_m4_i0_i0 (.D(n2285[0]), .SP(clk_N_683_enable_392), .CD(n14361), 
            .CK(clk_N_683), .Q(PWMdut_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i0.GSR = "DISABLED";
    LUT4 i13360_2_lut (.A(addOut[10]), .B(n22105), .Z(backOut3_28__N_1678[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13360_2_lut.init = 16'h2222;
    LUT4 mux_1241_i12_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[11]), 
         .D(speed_set_m4[11]), .Z(n2581[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i12_3_lut_4_lut.init = 16'hfe10;
    FD1P3IX dutyout_m3_i0_i0 (.D(n2273[0]), .SP(clk_N_683_enable_392), .CD(n14352), 
            .CK(clk_N_683), .Q(PWMdut_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i0.GSR = "DISABLED";
    FD1P3IX intgOut1_i0 (.D(addOut[0]), .SP(clk_N_683_enable_390), .CD(n14250), 
            .CK(clk_N_683), .Q(intgOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i0.GSR = "ENABLED";
    LUT4 i2_4_lut_then_3_lut_adj_124 (.A(ss[2]), .B(n22105), .C(ss[1]), 
         .Z(n21392)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_4_lut_then_3_lut_adj_124.init = 16'hfefe;
    CCU2D addOut_2081_add_4_15 (.A0(multOut[13]), .B0(n16396), .C0(addOut[13]), 
          .D0(addIn2_28__N_1246[13]), .A1(multOut[14]), .B1(n16396), .C1(addOut[14]), 
          .D1(addIn2_28__N_1246[14]), .CIN(n18224), .COUT(n18225), .S0(n121[13]), 
          .S1(n121[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_15.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_15.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_15.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_15.INJECT1_1 = "NO";
    CCU2D add_14998_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18391), 
          .S0(n3720));
    defparam add_14998_cout.INIT0 = 16'h0000;
    defparam add_14998_cout.INIT1 = 16'h0000;
    defparam add_14998_cout.INJECT1_0 = "NO";
    defparam add_14998_cout.INJECT1_1 = "NO";
    FD1P3IX dutyout_m2_i0_i0 (.D(n2261[0]), .SP(clk_N_683_enable_392), .CD(n14343), 
            .CK(clk_N_683), .Q(PWMdut_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i0.GSR = "DISABLED";
    LUT4 i13359_2_lut (.A(addOut[9]), .B(n22105), .Z(backOut3_28__N_1678[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13359_2_lut.init = 16'h2222;
    LUT4 i2_3_lut_4_lut_adj_125 (.A(n21298), .B(n21297), .C(n21317), .D(n21299), 
         .Z(n7_c)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i2_3_lut_4_lut_adj_125.init = 16'hffef;
    LUT4 mux_1241_i13_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[12]), 
         .D(speed_set_m4[12]), .Z(n2581[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13674_2_lut_rep_313 (.A(n15694), .B(n49), .Z(n21294)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13674_2_lut_rep_313.init = 16'heeee;
    PFUMX mux_137_i29 (.BLUT(n581[28]), .ALUT(intgOut3[28]), .C0(n21308), 
          .Z(n611[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    CCU2D add_14998_20 (.A0(speed_set_m3[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18390), .COUT(n18391));
    defparam add_14998_20.INIT0 = 16'h5aaa;
    defparam add_14998_20.INIT1 = 16'h0aaa;
    defparam add_14998_20.INJECT1_0 = "NO";
    defparam add_14998_20.INJECT1_1 = "NO";
    CCU2D add_14998_18 (.A0(speed_set_m3[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18389), .COUT(n18390));
    defparam add_14998_18.INIT0 = 16'h5aaa;
    defparam add_14998_18.INIT1 = 16'h5aaa;
    defparam add_14998_18.INJECT1_0 = "NO";
    defparam add_14998_18.INJECT1_1 = "NO";
    CCU2D add_1172_7 (.A0(n1328[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1328[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18142), 
          .COUT(n18143), .S0(n2273[5]), .S1(n2273[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1172_7.INIT0 = 16'hf555;
    defparam add_1172_7.INIT1 = 16'hf555;
    defparam add_1172_7.INJECT1_0 = "NO";
    defparam add_1172_7.INJECT1_1 = "NO";
    LUT4 i11709_3_lut_4_lut (.A(n1061), .B(n3832), .C(n21311), .D(clk_N_683_enable_331), 
         .Z(n14278)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i11709_3_lut_4_lut.init = 16'hfe00;
    LUT4 i13358_2_lut (.A(addOut[8]), .B(n22105), .Z(backOut3_28__N_1678[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13358_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_else_3_lut (.A(ss[2]), .B(n22105), .C(ss[1]), .D(ss[3]), 
         .Z(n21391)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i2_4_lut_else_3_lut.init = 16'hffef;
    LUT4 i3_2_lut_adj_126 (.A(speed_set_m1[18]), .B(speed_set_m1[5]), .Z(n24_adj_2193)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i3_2_lut_adj_126.init = 16'heeee;
    CCU2D addOut_2081_add_4_13 (.A0(multOut[11]), .B0(n16396), .C0(addOut[11]), 
          .D0(addIn2_28__N_1246[11]), .A1(multOut[12]), .B1(n16396), .C1(addOut[12]), 
          .D1(addIn2_28__N_1246[12]), .CIN(n18223), .COUT(n18224), .S0(n121[11]), 
          .S1(n121[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_13.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_13.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_13.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_13.INJECT1_1 = "NO";
    LUT4 i13355_2_lut (.A(addOut[7]), .B(n22105), .Z(backOut3_28__N_1678[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13355_2_lut.init = 16'h2222;
    LUT4 mux_1241_i15_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[14]), 
         .D(speed_set_m4[14]), .Z(n2581[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_91_i13_3_lut_4_lut_4_lut (.A(n21308), .B(\speed_avg_m4[12] ), 
         .C(n4322), .D(n22082), .Z(n367[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i13_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_1241_i16_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[15]), 
         .D(speed_set_m4[15]), .Z(n2581[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13143_2_lut_rep_405 (.A(ss[0]), .B(ss[1]), .Z(n22083)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13143_2_lut_rep_405.init = 16'h8888;
    LUT4 i2_4_lut_else_3_lut_4_lut (.A(n22105), .B(ss[0]), .C(ss[1]), 
         .D(ss[2]), .Z(n21388)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(C (D)))) */ ;
    defparam i2_4_lut_else_3_lut_4_lut.init = 16'hebff;
    LUT4 mux_1241_i2_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[1]), 
         .D(speed_set_m4[1]), .Z(n2581[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i2_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_14998_16 (.A0(speed_set_m3[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18388), .COUT(n18389));
    defparam add_14998_16.INIT0 = 16'h5aaa;
    defparam add_14998_16.INIT1 = 16'h5aaa;
    defparam add_14998_16.INJECT1_0 = "NO";
    defparam add_14998_16.INJECT1_1 = "NO";
    FD1P3IX dutyout_m1_i0_i0 (.D(n2249[0]), .SP(clk_N_683_enable_392), .CD(n14334), 
            .CK(clk_N_683), .Q(PWMdut_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i0.GSR = "DISABLED";
    LUT4 i2_4_lut_then_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(ss[2]), .D(n22105), 
         .Z(n21389)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_4_lut_then_3_lut_4_lut.init = 16'hfff7;
    LUT4 mux_91_i10_3_lut_4_lut_4_lut (.A(n21308), .B(\speed_avg_m4[9] ), 
         .C(n4322), .D(n22082), .Z(n367[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i10_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 i2_4_lut_else_3_lut_adj_127 (.A(ss[0]), .B(ss[2]), .C(n22084), 
         .D(n21325), .Z(n22093)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;
    defparam i2_4_lut_else_3_lut_adj_127.init = 16'hfb00;
    LUT4 i1_4_lut_then_4_lut (.A(n22105), .B(ss[0]), .C(ss[1]), .D(ss[3]), 
         .Z(n21398)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_else_4_lut (.A(n22105), .B(ss[0]), .C(ss[1]), .D(ss[3]), 
         .Z(n21397)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0100;
    LUT4 i13114_2_lut_rep_406 (.A(n22105), .B(ss[3]), .Z(n22084)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13114_2_lut_rep_406.init = 16'heeee;
    LUT4 i17139_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut (.A(n22105), .B(ss[3]), 
         .C(n4328), .D(n21359), .Z(n20272)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i17139_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 mux_91_i9_3_lut_4_lut_4_lut (.A(n21308), .B(\speed_avg_m4[8] ), 
         .C(n4322), .D(n22082), .Z(n367[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i9_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_1241_i17_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[16]), 
         .D(speed_set_m4[16]), .Z(n2581[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i17_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_189_i18_3_lut_3_lut (.A(n1061), .B(n3832), .C(addOut[17]), 
         .Z(intgOut0_28__N_1433[17])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i18_3_lut_3_lut.init = 16'hbaba;
    LUT4 i13352_2_lut (.A(addOut[6]), .B(n22105), .Z(backOut3_28__N_1678[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13352_2_lut.init = 16'h2222;
    LUT4 mux_1241_i18_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[17]), 
         .D(speed_set_m4[17]), .Z(n2581[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i18_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i20_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[19]), 
         .D(speed_set_m4[19]), .Z(n2581[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i20_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i21_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[20]), 
         .D(speed_set_m4[20]), .Z(n2581[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i14_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[13]), 
         .D(speed_set_m4[13]), .Z(n2581[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i14_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_189_i17_3_lut_3_lut (.A(n1061), .B(n3832), .C(addOut[16]), 
         .Z(intgOut0_28__N_1433[16])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i17_3_lut_3_lut.init = 16'hbaba;
    CCU2D add_14998_14 (.A0(speed_set_m3[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18387), .COUT(n18388));
    defparam add_14998_14.INIT0 = 16'h5555;
    defparam add_14998_14.INIT1 = 16'h5aaa;
    defparam add_14998_14.INJECT1_0 = "NO";
    defparam add_14998_14.INJECT1_1 = "NO";
    CCU2D add_1172_5 (.A0(n1328[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1328[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18141), 
          .COUT(n18142), .S0(n2273[3]), .S1(n2273[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1172_5.INIT0 = 16'hf555;
    defparam add_1172_5.INIT1 = 16'hf555;
    defparam add_1172_5.INJECT1_0 = "NO";
    defparam add_1172_5.INJECT1_1 = "NO";
    CCU2D add_1172_3 (.A0(n1328[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1328[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18140), 
          .COUT(n18141), .S0(n2273[1]), .S1(n2273[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1172_3.INIT0 = 16'hf555;
    defparam add_1172_3.INIT1 = 16'hf555;
    defparam add_1172_3.INJECT1_0 = "NO";
    defparam add_1172_3.INJECT1_1 = "NO";
    CCU2D add_14998_12 (.A0(speed_set_m3[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18386), .COUT(n18387));
    defparam add_14998_12.INIT0 = 16'h5aaa;
    defparam add_14998_12.INIT1 = 16'h5aaa;
    defparam add_14998_12.INJECT1_0 = "NO";
    defparam add_14998_12.INJECT1_1 = "NO";
    CCU2D add_14998_10 (.A0(speed_set_m3[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18385), .COUT(n18386));
    defparam add_14998_10.INIT0 = 16'h5555;
    defparam add_14998_10.INIT1 = 16'h5555;
    defparam add_14998_10.INJECT1_0 = "NO";
    defparam add_14998_10.INJECT1_1 = "NO";
    PFUMX mux_137_i1 (.BLUT(n581[0]), .ALUT(intgOut3[0]), .C0(n21308), 
          .Z(n611[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=311, LSE_RLINE=311 */ ;
    LUT4 mux_189_i15_3_lut_3_lut (.A(n1061), .B(n3832), .C(addOut[14]), 
         .Z(intgOut0_28__N_1433[14])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i15_3_lut_3_lut.init = 16'hbaba;
    LUT4 mux_1241_i3_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[2]), 
         .D(speed_set_m4[2]), .Z(n2581[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i3_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1172_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1328[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18140), 
          .S1(n2273[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1172_1.INIT0 = 16'hF000;
    defparam add_1172_1.INIT1 = 16'h0aaa;
    defparam add_1172_1.INJECT1_0 = "NO";
    defparam add_1172_1.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_11 (.A0(multOut[9]), .B0(n16396), .C0(addOut[9]), 
          .D0(addIn2_28__N_1246[9]), .A1(multOut[10]), .B1(n16396), .C1(addOut[10]), 
          .D1(addIn2_28__N_1246[10]), .CIN(n18222), .COUT(n18223), .S0(n121[9]), 
          .S1(n121[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_11.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_11.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_11.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_11.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_9 (.A0(multOut[7]), .B0(n16396), .C0(addOut[7]), 
          .D0(addIn2_28__N_1246[7]), .A1(multOut[8]), .B1(n16396), .C1(addOut[8]), 
          .D1(addIn2_28__N_1246[8]), .CIN(n18221), .COUT(n18222), .S0(n121[7]), 
          .S1(n121[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_9.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_9.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_9.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_9.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_7 (.A0(multOut[5]), .B0(n16396), .C0(addOut[5]), 
          .D0(addIn2_28__N_1246[5]), .A1(multOut[6]), .B1(n16396), .C1(addOut[6]), 
          .D1(addIn2_28__N_1246[6]), .CIN(n18220), .COUT(n18221), .S0(n121[5]), 
          .S1(n121[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_7.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_7.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_7.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_7.INJECT1_1 = "NO";
    CCU2D add_1171_11 (.A0(n1307[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18139), 
          .S0(n2261[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1171_11.INIT0 = 16'hf555;
    defparam add_1171_11.INIT1 = 16'h0000;
    defparam add_1171_11.INJECT1_0 = "NO";
    defparam add_1171_11.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_5 (.A0(multOut[3]), .B0(n16396), .C0(addOut[3]), 
          .D0(addIn2_28__N_1246[3]), .A1(multOut[4]), .B1(n16396), .C1(addOut[4]), 
          .D1(addIn2_28__N_1246[4]), .CIN(n18219), .COUT(n18220), .S0(n121[3]), 
          .S1(n121[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_5.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_5.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_5.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_5.INJECT1_1 = "NO";
    CCU2D add_14998_8 (.A0(speed_set_m3[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18384), .COUT(n18385));
    defparam add_14998_8.INIT0 = 16'h5aaa;
    defparam add_14998_8.INIT1 = 16'h5555;
    defparam add_14998_8.INJECT1_0 = "NO";
    defparam add_14998_8.INJECT1_1 = "NO";
    CCU2D add_1171_9 (.A0(n1307[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1307[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18138), 
          .COUT(n18139), .S0(n2261[7]), .S1(n2261[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1171_9.INIT0 = 16'hf555;
    defparam add_1171_9.INIT1 = 16'hf555;
    defparam add_1171_9.INJECT1_0 = "NO";
    defparam add_1171_9.INJECT1_1 = "NO";
    CCU2D add_1171_7 (.A0(n1307[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1307[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18137), 
          .COUT(n18138), .S0(n2261[5]), .S1(n2261[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1171_7.INIT0 = 16'hf555;
    defparam add_1171_7.INIT1 = 16'hf555;
    defparam add_1171_7.INJECT1_0 = "NO";
    defparam add_1171_7.INJECT1_1 = "NO";
    LUT4 mux_189_i10_3_lut_3_lut (.A(n1061), .B(n3832), .C(addOut[9]), 
         .Z(intgOut0_28__N_1433[9])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i10_3_lut_3_lut.init = 16'hbaba;
    CCU2D add_14998_6 (.A0(speed_set_m3[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18383), .COUT(n18384));
    defparam add_14998_6.INIT0 = 16'h5aaa;
    defparam add_14998_6.INIT1 = 16'h5aaa;
    defparam add_14998_6.INJECT1_0 = "NO";
    defparam add_14998_6.INJECT1_1 = "NO";
    CCU2D add_14998_4 (.A0(speed_set_m3[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18382), .COUT(n18383));
    defparam add_14998_4.INIT0 = 16'h5555;
    defparam add_14998_4.INIT1 = 16'h5aaa;
    defparam add_14998_4.INJECT1_0 = "NO";
    defparam add_14998_4.INJECT1_1 = "NO";
    CCU2D add_14998_2 (.A0(speed_set_m3[1]), .B0(speed_set_m3[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18382));
    defparam add_14998_2.INIT0 = 16'h1000;
    defparam add_14998_2.INIT1 = 16'h5555;
    defparam add_14998_2.INJECT1_0 = "NO";
    defparam add_14998_2.INJECT1_1 = "NO";
    CCU2D add_14999_17 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18381), .S1(n3696));
    defparam add_14999_17.INIT0 = 16'h5555;
    defparam add_14999_17.INIT1 = 16'h0000;
    defparam add_14999_17.INJECT1_0 = "NO";
    defparam add_14999_17.INJECT1_1 = "NO";
    CCU2D add_14999_15 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18380), .COUT(n18381));
    defparam add_14999_15.INIT0 = 16'hf555;
    defparam add_14999_15.INIT1 = 16'hf555;
    defparam add_14999_15.INJECT1_0 = "NO";
    defparam add_14999_15.INJECT1_1 = "NO";
    CCU2D add_14999_13 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18379), .COUT(n18380));
    defparam add_14999_13.INIT0 = 16'hf555;
    defparam add_14999_13.INIT1 = 16'hf555;
    defparam add_14999_13.INJECT1_0 = "NO";
    defparam add_14999_13.INJECT1_1 = "NO";
    CCU2D add_14999_11 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18378), .COUT(n18379));
    defparam add_14999_11.INIT0 = 16'hf555;
    defparam add_14999_11.INIT1 = 16'hf555;
    defparam add_14999_11.INJECT1_0 = "NO";
    defparam add_14999_11.INJECT1_1 = "NO";
    CCU2D add_14999_9 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18377), .COUT(n18378));
    defparam add_14999_9.INIT0 = 16'hf555;
    defparam add_14999_9.INIT1 = 16'h0aaa;
    defparam add_14999_9.INJECT1_0 = "NO";
    defparam add_14999_9.INJECT1_1 = "NO";
    CCU2D add_14999_7 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18376), .COUT(n18377));
    defparam add_14999_7.INIT0 = 16'h0aaa;
    defparam add_14999_7.INIT1 = 16'hf555;
    defparam add_14999_7.INJECT1_0 = "NO";
    defparam add_14999_7.INJECT1_1 = "NO";
    CCU2D add_14999_5 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18375), .COUT(n18376));
    defparam add_14999_5.INIT0 = 16'h0aaa;
    defparam add_14999_5.INIT1 = 16'h0aaa;
    defparam add_14999_5.INJECT1_0 = "NO";
    defparam add_14999_5.INJECT1_1 = "NO";
    CCU2D add_14999_3 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18374), .COUT(n18375));
    defparam add_14999_3.INIT0 = 16'hf555;
    defparam add_14999_3.INIT1 = 16'hf555;
    defparam add_14999_3.INJECT1_0 = "NO";
    defparam add_14999_3.INJECT1_1 = "NO";
    CCU2D add_14999_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[4]), .B1(speed_set_m3[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18374));
    defparam add_14999_1.INIT0 = 16'hF000;
    defparam add_14999_1.INIT1 = 16'ha666;
    defparam add_14999_1.INJECT1_0 = "NO";
    defparam add_14999_1.INJECT1_1 = "NO";
    CCU2D add_15000_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18373), 
          .S0(n3672));
    defparam add_15000_cout.INIT0 = 16'h0000;
    defparam add_15000_cout.INIT1 = 16'h0000;
    defparam add_15000_cout.INJECT1_0 = "NO";
    defparam add_15000_cout.INJECT1_1 = "NO";
    CCU2D add_15000_20 (.A0(speed_set_m2[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18372), .COUT(n18373));
    defparam add_15000_20.INIT0 = 16'h5aaa;
    defparam add_15000_20.INIT1 = 16'h0aaa;
    defparam add_15000_20.INJECT1_0 = "NO";
    defparam add_15000_20.INJECT1_1 = "NO";
    CCU2D add_15000_18 (.A0(speed_set_m2[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18371), .COUT(n18372));
    defparam add_15000_18.INIT0 = 16'h5aaa;
    defparam add_15000_18.INIT1 = 16'h5aaa;
    defparam add_15000_18.INJECT1_0 = "NO";
    defparam add_15000_18.INJECT1_1 = "NO";
    CCU2D add_15000_16 (.A0(speed_set_m2[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18370), .COUT(n18371));
    defparam add_15000_16.INIT0 = 16'h5aaa;
    defparam add_15000_16.INIT1 = 16'h5aaa;
    defparam add_15000_16.INJECT1_0 = "NO";
    defparam add_15000_16.INJECT1_1 = "NO";
    CCU2D add_15000_14 (.A0(speed_set_m2[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18369), .COUT(n18370));
    defparam add_15000_14.INIT0 = 16'h5555;
    defparam add_15000_14.INIT1 = 16'h5aaa;
    defparam add_15000_14.INJECT1_0 = "NO";
    defparam add_15000_14.INJECT1_1 = "NO";
    CCU2D add_15000_12 (.A0(speed_set_m2[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18368), .COUT(n18369));
    defparam add_15000_12.INIT0 = 16'h5aaa;
    defparam add_15000_12.INIT1 = 16'h5aaa;
    defparam add_15000_12.INJECT1_0 = "NO";
    defparam add_15000_12.INJECT1_1 = "NO";
    CCU2D add_15000_10 (.A0(speed_set_m2[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18367), .COUT(n18368));
    defparam add_15000_10.INIT0 = 16'h5555;
    defparam add_15000_10.INIT1 = 16'h5555;
    defparam add_15000_10.INJECT1_0 = "NO";
    defparam add_15000_10.INJECT1_1 = "NO";
    CCU2D add_15000_8 (.A0(speed_set_m2[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18366), .COUT(n18367));
    defparam add_15000_8.INIT0 = 16'h5aaa;
    defparam add_15000_8.INIT1 = 16'h5555;
    defparam add_15000_8.INJECT1_0 = "NO";
    defparam add_15000_8.INJECT1_1 = "NO";
    CCU2D add_15000_6 (.A0(speed_set_m2[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18365), .COUT(n18366));
    defparam add_15000_6.INIT0 = 16'h5aaa;
    defparam add_15000_6.INIT1 = 16'h5aaa;
    defparam add_15000_6.INJECT1_0 = "NO";
    defparam add_15000_6.INJECT1_1 = "NO";
    CCU2D add_15000_4 (.A0(speed_set_m2[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18364), .COUT(n18365));
    defparam add_15000_4.INIT0 = 16'h5555;
    defparam add_15000_4.INIT1 = 16'h5aaa;
    defparam add_15000_4.INJECT1_0 = "NO";
    defparam add_15000_4.INJECT1_1 = "NO";
    PFUMX i17321 (.BLUT(n21397), .ALUT(n21398), .C0(ss[2]), .Z(n4322));
    CCU2D add_223_17 (.A0(Out3[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18064), 
          .S0(n1349[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_17.INIT0 = 16'h5aaa;
    defparam add_223_17.INIT1 = 16'h0000;
    defparam add_223_17.INJECT1_0 = "NO";
    defparam add_223_17.INJECT1_1 = "NO";
    CCU2D add_223_15 (.A0(Out3[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18063), 
          .COUT(n18064), .S0(n1349[13]), .S1(n1349[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_15.INIT0 = 16'h5aaa;
    defparam add_223_15.INIT1 = 16'h5aaa;
    defparam add_223_15.INJECT1_0 = "NO";
    defparam add_223_15.INJECT1_1 = "NO";
    CCU2D add_223_13 (.A0(Out3[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18062), 
          .COUT(n18063), .S0(n1349[11]), .S1(n1349[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_13.INIT0 = 16'h5aaa;
    defparam add_223_13.INIT1 = 16'h5aaa;
    defparam add_223_13.INJECT1_0 = "NO";
    defparam add_223_13.INJECT1_1 = "NO";
    CCU2D add_223_11 (.A0(Out3[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18061), 
          .COUT(n18062), .S0(n1349[9]), .S1(n1349[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_11.INIT0 = 16'h5aaa;
    defparam add_223_11.INIT1 = 16'h5aaa;
    defparam add_223_11.INJECT1_0 = "NO";
    defparam add_223_11.INJECT1_1 = "NO";
    CCU2D add_1171_5 (.A0(n1307[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1307[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18136), 
          .COUT(n18137), .S0(n2261[3]), .S1(n2261[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1171_5.INIT0 = 16'hf555;
    defparam add_1171_5.INIT1 = 16'hf555;
    defparam add_1171_5.INJECT1_0 = "NO";
    defparam add_1171_5.INJECT1_1 = "NO";
    CCU2D add_1171_3 (.A0(n1307[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1307[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18135), 
          .COUT(n18136), .S0(n2261[1]), .S1(n2261[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1171_3.INIT0 = 16'hf555;
    defparam add_1171_3.INIT1 = 16'hf555;
    defparam add_1171_3.INJECT1_0 = "NO";
    defparam add_1171_3.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_3 (.A0(multOut[1]), .B0(n16396), .C0(addOut[1]), 
          .D0(addIn2_28__N_1246[1]), .A1(multOut[2]), .B1(n16396), .C1(addOut[2]), 
          .D1(addIn2_28__N_1246[2]), .CIN(n18218), .COUT(n18219), .S0(n121[1]), 
          .S1(n121[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_3.INIT0 = 16'h569a;
    defparam addOut_2081_add_4_3.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_3.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_3.INJECT1_1 = "NO";
    CCU2D add_15000_2 (.A0(speed_set_m2[1]), .B0(speed_set_m2[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18364));
    defparam add_15000_2.INIT0 = 16'h1000;
    defparam add_15000_2.INIT1 = 16'h5555;
    defparam add_15000_2.INJECT1_0 = "NO";
    defparam add_15000_2.INJECT1_1 = "NO";
    CCU2D add_15001_17 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18363), .S1(n3648));
    defparam add_15001_17.INIT0 = 16'h5555;
    defparam add_15001_17.INIT1 = 16'h0000;
    defparam add_15001_17.INJECT1_0 = "NO";
    defparam add_15001_17.INJECT1_1 = "NO";
    CCU2D add_223_9 (.A0(Out3[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18060), 
          .COUT(n18061), .S0(n1349[7]), .S1(n1349[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_9.INIT0 = 16'h5aaa;
    defparam add_223_9.INIT1 = 16'h5aaa;
    defparam add_223_9.INJECT1_0 = "NO";
    defparam add_223_9.INJECT1_1 = "NO";
    CCU2D add_223_7 (.A0(Out3[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18059), 
          .COUT(n18060), .S0(n1349[5]), .S1(n1349[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_7.INIT0 = 16'h5aaa;
    defparam add_223_7.INIT1 = 16'h5aaa;
    defparam add_223_7.INJECT1_0 = "NO";
    defparam add_223_7.INJECT1_1 = "NO";
    CCU2D add_223_5 (.A0(Out3[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18058), 
          .COUT(n18059), .S0(n1349[3]), .S1(n1349[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_5.INIT0 = 16'h5aaa;
    defparam add_223_5.INIT1 = 16'h5aaa;
    defparam add_223_5.INJECT1_0 = "NO";
    defparam add_223_5.INJECT1_1 = "NO";
    CCU2D add_223_3 (.A0(Out3[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18057), 
          .COUT(n18058), .S0(n1349[1]), .S1(n1349[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_3.INIT0 = 16'h5aaa;
    defparam add_223_3.INIT1 = 16'h5aaa;
    defparam add_223_3.INJECT1_0 = "NO";
    defparam add_223_3.INJECT1_1 = "NO";
    CCU2D add_1171_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1307[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18135), 
          .S1(n2261[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1171_1.INIT0 = 16'hF000;
    defparam add_1171_1.INIT1 = 16'h0aaa;
    defparam add_1171_1.INJECT1_0 = "NO";
    defparam add_1171_1.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_23 (.A0(n2341[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2341[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18133), .S0(n4415), .S1(n4414));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_23.INIT0 = 16'h5555;
    defparam sub_16_rep_3_add_2_23.INIT1 = 16'h5555;
    defparam sub_16_rep_3_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_23.INJECT1_1 = "NO";
    CCU2D addOut_2081_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(multOut[0]), .B1(n16396), .C1(addOut[0]), 
          .D1(addIn2_28__N_1246[0]), .COUT(n18218), .S1(n121[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081_add_4_1.INIT0 = 16'hF000;
    defparam addOut_2081_add_4_1.INIT1 = 16'h569a;
    defparam addOut_2081_add_4_1.INJECT1_0 = "NO";
    defparam addOut_2081_add_4_1.INJECT1_1 = "NO";
    CCU2D add_15001_15 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18362), .COUT(n18363));
    defparam add_15001_15.INIT0 = 16'hf555;
    defparam add_15001_15.INIT1 = 16'hf555;
    defparam add_15001_15.INJECT1_0 = "NO";
    defparam add_15001_15.INJECT1_1 = "NO";
    CCU2D add_15001_13 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18361), .COUT(n18362));
    defparam add_15001_13.INIT0 = 16'hf555;
    defparam add_15001_13.INIT1 = 16'hf555;
    defparam add_15001_13.INJECT1_0 = "NO";
    defparam add_15001_13.INJECT1_1 = "NO";
    PFUMX i17317 (.BLUT(n21391), .ALUT(n21392), .C0(ss[0]), .Z(n16470));
    FD1S3AX addOut_2081__i1 (.D(n121[1]), .CK(clk_N_683), .Q(addOut[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i1.GSR = "ENABLED";
    LUT4 i13225_2_lut_3_lut (.A(n1061), .B(n3832), .C(addOut[6]), .Z(intgOut0_28__N_1433[6])) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i13225_2_lut_3_lut.init = 16'hfefe;
    LUT4 i11681_3_lut_4_lut (.A(n1061), .B(n3832), .C(n21313), .D(clk_N_683_enable_390), 
         .Z(n14250)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i11681_3_lut_4_lut.init = 16'hfe00;
    LUT4 i13676_2_lut_rep_314_4_lut (.A(n9_adj_2138), .B(n9_adj_2137), .C(n21326), 
         .D(n56), .Z(n21295)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i13676_2_lut_rep_314_4_lut.init = 16'hff80;
    LUT4 mux_1241_i4_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[3]), 
         .D(speed_set_m4[3]), .Z(n2581[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i8_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[7]), 
         .D(speed_set_m4[7]), .Z(n2581[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i1_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[0]), 
         .D(speed_set_m4[0]), .Z(n2581[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i7_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[6]), 
         .D(speed_set_m4[6]), .Z(n2581[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1241_i9_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[8]), 
         .D(speed_set_m4[8]), .Z(n2581[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i9_3_lut_4_lut.init = 16'hfe10;
    PFUMX i17315 (.BLUT(n21388), .ALUT(n21389), .C0(ss[3]), .Z(n15694));
    LUT4 i17102_4_lut_4_lut (.A(n21325), .B(n20022), .C(n21326), .D(n21320), 
         .Z(n20045)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 185[26])
    defparam i17102_4_lut_4_lut.init = 16'hdfff;
    LUT4 mux_1241_i10_3_lut_4_lut (.A(n15694), .B(n49), .C(speed_set_m3[9]), 
         .D(speed_set_m4[9]), .Z(n2581[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1241_i10_3_lut_4_lut.init = 16'hfe10;
    FD1S3AX addOut_2081__i2 (.D(n121[2]), .CK(clk_N_683), .Q(addOut[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i2.GSR = "ENABLED";
    FD1S3AX addOut_2081__i3 (.D(n121[3]), .CK(clk_N_683), .Q(addOut[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i3.GSR = "ENABLED";
    FD1S3AX addOut_2081__i4 (.D(n121[4]), .CK(clk_N_683), .Q(addOut[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i4.GSR = "ENABLED";
    FD1S3AX addOut_2081__i5 (.D(n121[5]), .CK(clk_N_683), .Q(addOut[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i5.GSR = "ENABLED";
    FD1S3AX addOut_2081__i6 (.D(n121[6]), .CK(clk_N_683), .Q(addOut[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i6.GSR = "ENABLED";
    FD1S3AX addOut_2081__i7 (.D(n121[7]), .CK(clk_N_683), .Q(addOut[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i7.GSR = "ENABLED";
    FD1S3AX addOut_2081__i8 (.D(n121[8]), .CK(clk_N_683), .Q(addOut[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i8.GSR = "ENABLED";
    FD1S3AX addOut_2081__i9 (.D(n121[9]), .CK(clk_N_683), .Q(addOut[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i9.GSR = "ENABLED";
    FD1S3AX addOut_2081__i10 (.D(n121[10]), .CK(clk_N_683), .Q(addOut[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i10.GSR = "ENABLED";
    FD1S3AX addOut_2081__i11 (.D(n121[11]), .CK(clk_N_683), .Q(addOut[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i11.GSR = "ENABLED";
    FD1S3AX addOut_2081__i12 (.D(n121[12]), .CK(clk_N_683), .Q(addOut[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i12.GSR = "ENABLED";
    FD1S3AX addOut_2081__i13 (.D(n121[13]), .CK(clk_N_683), .Q(addOut[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i13.GSR = "ENABLED";
    FD1S3AX addOut_2081__i14 (.D(n121[14]), .CK(clk_N_683), .Q(addOut[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i14.GSR = "ENABLED";
    FD1S3AX addOut_2081__i15 (.D(n121[15]), .CK(clk_N_683), .Q(addOut[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i15.GSR = "ENABLED";
    FD1S3AX addOut_2081__i16 (.D(n121[16]), .CK(clk_N_683), .Q(addOut[16])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i16.GSR = "ENABLED";
    FD1S3AX addOut_2081__i17 (.D(n121[17]), .CK(clk_N_683), .Q(addOut[17])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i17.GSR = "ENABLED";
    FD1S3AX addOut_2081__i18 (.D(n121[18]), .CK(clk_N_683), .Q(addOut[18])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i18.GSR = "ENABLED";
    FD1S3AX addOut_2081__i19 (.D(n121[19]), .CK(clk_N_683), .Q(addOut[19])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i19.GSR = "ENABLED";
    FD1S3AX addOut_2081__i20 (.D(n121[20]), .CK(clk_N_683), .Q(addOut[20])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i20.GSR = "ENABLED";
    FD1S3AX addOut_2081__i21 (.D(n121[21]), .CK(clk_N_683), .Q(addOut[21])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i21.GSR = "ENABLED";
    FD1S3AX addOut_2081__i22 (.D(n121[22]), .CK(clk_N_683), .Q(addOut[22])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i22.GSR = "ENABLED";
    FD1S3AX addOut_2081__i23 (.D(n121[23]), .CK(clk_N_683), .Q(addOut[23])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i23.GSR = "ENABLED";
    FD1S3AX addOut_2081__i24 (.D(n121[24]), .CK(clk_N_683), .Q(addOut[24])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i24.GSR = "ENABLED";
    FD1S3AX addOut_2081__i25 (.D(n121[25]), .CK(clk_N_683), .Q(addOut[25])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i25.GSR = "ENABLED";
    FD1S3AX addOut_2081__i26 (.D(n121[26]), .CK(clk_N_683), .Q(addOut[26])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i26.GSR = "ENABLED";
    FD1S3AX addOut_2081__i27 (.D(n121[27]), .CK(clk_N_683), .Q(addOut[27])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i27.GSR = "ENABLED";
    FD1S3AX addOut_2081__i28 (.D(n121[28]), .CK(clk_N_683), .Q(addOut[28])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2081__i28.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module HALL_U5
//

module HALL_U5 (clk_1mhz, n22097, \speed_m1[0] , hallsense_m1, rst, 
            clkout_c_enable_173, H_A_m1_c, H_B_m1_c, H_C_m1_c, \speed_m1[1] , 
            \speed_m1[2] , \speed_m1[3] , \speed_m1[4] , \speed_m1[5] , 
            \speed_m1[6] , \speed_m1[7] , \speed_m1[8] , \speed_m1[9] , 
            \speed_m1[10] , \speed_m1[11] , \speed_m1[12] , \speed_m1[13] , 
            \speed_m1[14] , \speed_m1[15] , \speed_m1[16] , \speed_m1[17] , 
            \speed_m1[18] , \speed_m1[19] , GND_net);
    input clk_1mhz;
    input n22097;
    output \speed_m1[0] ;
    output [2:0]hallsense_m1;
    input rst;
    input clkout_c_enable_173;
    input H_A_m1_c;
    input H_B_m1_c;
    input H_C_m1_c;
    output \speed_m1[1] ;
    output \speed_m1[2] ;
    output \speed_m1[3] ;
    output \speed_m1[4] ;
    output \speed_m1[5] ;
    output \speed_m1[6] ;
    output \speed_m1[7] ;
    output \speed_m1[8] ;
    output \speed_m1[9] ;
    output \speed_m1[10] ;
    output \speed_m1[11] ;
    output \speed_m1[12] ;
    output \speed_m1[13] ;
    output \speed_m1[14] ;
    output \speed_m1[15] ;
    output \speed_m1[16] ;
    output \speed_m1[17] ;
    output \speed_m1[18] ;
    output \speed_m1[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_63;
    wire [19:0]count_19__N_1873;
    
    wire stable_counting, clk_1mhz_enable_3, n14400;
    wire [19:0]speedt_19__N_1853;
    
    wire hall3_lat, n11414, n11427, stable_counting_N_1935, n19413, 
        n19584, n19790, n19738;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4545;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21338, n21303, n4, n19596, n19734, n21315, n19397, n19516, 
        hall3_old, n4_adj_2132, n21330;
    wire [6:0]n63;
    
    wire n21301, hall1_old, hall1_lat, hall2_old, hall2_lat, n12, 
        n21364, n21314, n21, n21322, n18082, n18081, n18080, n18079, 
        n18078, n18077, n18076, n18075, n18074, n18073, n18689, 
        n19634, n24, n20, n18;
    
    FD1P3AX speedt_i0_i0 (.D(count_19__N_1873[0]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22097), .SP(clk_1mhz_enable_3), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1853[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    LUT4 i11516_4_lut (.A(n11414), .B(n11427), .C(stable_counting), .D(stable_counting_N_1935), 
         .Z(clk_1mhz_enable_63)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11516_4_lut.init = 16'hcaea;
    LUT4 i1_4_lut (.A(n19413), .B(n19584), .C(n19790), .D(n19738), .Z(n11414)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0002;
    FD1S3IX count__i0 (.D(count_19__N_1873[0]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    LUT4 i2388_2_lut_rep_322_3_lut_4_lut (.A(stable_count[3]), .B(n21338), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21303)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2388_2_lut_rep_322_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21338), .C(stable_count[0]), 
         .D(stable_count[4]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h7f8f;
    LUT4 i16200_2_lut (.A(count[18]), .B(count[1]), .Z(n19584)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16200_2_lut.init = 16'heeee;
    LUT4 i16399_4_lut (.A(n19596), .B(n19734), .C(count[19]), .D(count[14]), 
         .Z(n19790)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16399_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut (.A(n21315), .B(stable_count[0]), .C(n19397), .D(n19516), 
         .Z(n11427)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_rep_349 (.A(hall3_old), .B(n4_adj_2132), .C(hall3_lat), 
         .Z(n21330)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_349.init = 16'hdede;
    LUT4 i2_4_lut (.A(n19516), .B(n63[2]), .C(n21301), .D(n4), .Z(stable_counting_N_1935)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i2_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4_adj_2132), .C(hall3_lat), 
         .D(n63[1]), .Z(n19516)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 i2360_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2360_2_lut.init = 16'h6666;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(rst), .CK(clk_1mhz), .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m1_c), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m1_c), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m1_c), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_1873[19]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_1873[18]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_1873[17]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_1873[16]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_1873[15]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_1873[14]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_1873[13]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_1873[12]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_1873[11]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_1873[10]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_1873[9]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_1873[8]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_1873[7]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_1873[6]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_1873[5]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_1873[4]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_1873[3]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_1873[2]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_1873[1]), .SP(clk_1mhz_enable_63), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    LUT4 i16212_2_lut (.A(count[17]), .B(count[12]), .Z(n19596)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16212_2_lut.init = 16'heeee;
    LUT4 i2238_2_lut (.A(stable_counting), .B(stable_counting_N_1935), .Z(n4545)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2238_2_lut.init = 16'h8888;
    FD1P3AX speed__i2 (.D(speedt_19__N_1853[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1853[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1853[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1853[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1853[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1853[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1853[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1853[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1853[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1853[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1853[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1853[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1853[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1853[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1853[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1853[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1853[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1853[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1853[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(count_19__N_1873[1]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_1873[2]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_1873[3]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_1873[4]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_1873[5]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_1873[6]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_1873[7]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_1873[8]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_1873[9]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_1873[10]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_1873[11]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_1873[12]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_1873[13]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_1873[14]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_1873[15]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_1873[16]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_1873[17]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_1873[18]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_1873[19]), .CK(clk_1mhz), .CD(n4545), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    LUT4 i6_4_lut (.A(count[2]), .B(n12), .C(count[9]), .D(count[8]), 
         .Z(n19413)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[3]), .B(count[10]), .C(count[13]), .D(count[0]), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i2383_2_lut_rep_333_3_lut_4_lut (.A(stable_count[2]), .B(n21364), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21314)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2383_2_lut_rep_333_3_lut_4_lut.init = 16'h8000;
    LUT4 i2381_2_lut_rep_334_3_lut_4_lut (.A(stable_count[2]), .B(n21364), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21315)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2381_2_lut_rep_334_3_lut_4_lut.init = 16'h78f0;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[0]), 
         .D(speedt[0]), .Z(speedt_19__N_1853[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[1]), 
         .D(speedt[1]), .Z(speedt_19__N_1853[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[2]), 
         .D(speedt[2]), .Z(speedt_19__N_1853[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[3]), 
         .D(speedt[3]), .Z(speedt_19__N_1853[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[4]), 
         .D(speedt[4]), .Z(speedt_19__N_1853[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[5]), 
         .D(speedt[5]), .Z(speedt_19__N_1853[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16345_3_lut_4_lut (.A(count[7]), .B(count[6]), .C(count[4]), 
         .D(count[11]), .Z(n19734)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16345_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[6]), 
         .D(speedt[6]), .Z(speedt_19__N_1853[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i8_2_lut_3_lut_4_lut (.A(count[5]), .B(count[16]), .C(count[6]), 
         .D(count[7]), .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i16349_2_lut_3_lut (.A(count[5]), .B(count[16]), .C(count[15]), 
         .Z(n19738)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16349_2_lut_3_lut.init = 16'hfefe;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[7]), 
         .D(speedt[7]), .Z(speedt_19__N_1853[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2362_2_lut_rep_383 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21364)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2362_2_lut_rep_383.init = 16'h8888;
    LUT4 i2367_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2367_2_lut_3_lut.init = 16'h7878;
    LUT4 i2369_2_lut_rep_357_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21338)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2369_2_lut_rep_357_3_lut.init = 16'h8080;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[8]), 
         .D(speedt[8]), .Z(speedt_19__N_1853[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[9]), 
         .D(speedt[9]), .Z(speedt_19__N_1853[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[10]), 
         .D(speedt[10]), .Z(speedt_19__N_1853[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2376_2_lut_rep_341_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21322)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2376_2_lut_rep_341_3_lut_4_lut.init = 16'h8000;
    LUT4 i2374_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2374_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[11]), 
         .D(speedt[11]), .Z(speedt_19__N_1853[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[12]), 
         .D(speedt[12]), .Z(speedt_19__N_1853[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[13]), 
         .D(speedt[13]), .Z(speedt_19__N_1853[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[14]), 
         .D(speedt[14]), .Z(speedt_19__N_1853[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[15]), 
         .D(speedt[15]), .Z(speedt_19__N_1853[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[16]), 
         .D(speedt[16]), .Z(speedt_19__N_1853[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[17]), 
         .D(speedt[17]), .Z(speedt_19__N_1853[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[18]), 
         .D(speedt[18]), .Z(speedt_19__N_1853[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11414), .B(n11427), .C(count_19__N_1873[19]), 
         .D(speedt[19]), .Z(speedt_19__N_1853[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21303), .SP(stable_counting), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21315), .SP(stable_counting), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18082), 
          .S0(count_19__N_1873[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18081), .COUT(n18082), .S0(count_19__N_1873[17]), .S1(count_19__N_1873[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18080), .COUT(n18081), .S0(count_19__N_1873[15]), .S1(count_19__N_1873[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18079), .COUT(n18080), .S0(count_19__N_1873[13]), .S1(count_19__N_1873[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18078), .COUT(n18079), .S0(count_19__N_1873[11]), .S1(count_19__N_1873[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18077), .COUT(n18078), .S0(count_19__N_1873[9]), .S1(count_19__N_1873[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18076), 
          .COUT(n18077), .S0(count_19__N_1873[7]), .S1(count_19__N_1873[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18075), 
          .COUT(n18076), .S0(count_19__N_1873[5]), .S1(count_19__N_1873[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_45 (.A(n21303), .B(n63[6]), .C(n63[3]), .D(n63[2]), 
         .Z(n19397)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_2_lut_4_lut_adj_45.init = 16'hfffe;
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18074), 
          .COUT(n18075), .S0(count_19__N_1873[3]), .S1(count_19__N_1873[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18073), 
          .COUT(n18074), .S0(count_19__N_1873[1]), .S1(count_19__N_1873[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14400), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=316, LSE_RLINE=316 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    LUT4 i2358_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2358_1_lut.init = 16'h5555;
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18073), 
          .S1(count_19__N_1873[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i17199_4_lut (.A(n18689), .B(n19634), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_3)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17199_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_46 (.A(n19596), .B(n19413), .C(n24), .D(n20), 
         .Z(n18689)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i1_4_lut_adj_46.init = 16'hfffb;
    LUT4 i2_3_lut_rep_320_4_lut (.A(stable_count[5]), .B(n21314), .C(n63[3]), 
         .D(n63[6]), .Z(n21301)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_320_4_lut.init = 16'hfff6;
    LUT4 i16249_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19634)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16249_4_lut.init = 16'h7bde;
    LUT4 i11_4_lut (.A(n21), .B(count[15]), .C(n18), .D(count[1]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut (.A(count[14]), .B(count[19]), .C(count[11]), .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i5_2_lut (.A(count[18]), .B(count[4]), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i11832_3_lut (.A(stable_counting), .B(n21330), .C(stable_counting_N_1935), 
         .Z(n14400)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i11832_3_lut.init = 16'ha8a8;
    LUT4 i2395_3_lut_4_lut (.A(stable_count[4]), .B(n21322), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2395_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_4_lut_adj_47 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4_adj_2132)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_47.init = 16'h7bde;
    
endmodule
//
// Verilog Description of module HALL_U3
//

module HALL_U3 (\speed_m3[0] , clk_1mhz, hallsense_m3, clkout_c_enable_173, 
            H_A_m3_c, H_B_m3_c, H_C_m3_c, rst, \speed_m3[1] , \speed_m3[2] , 
            \speed_m3[3] , \speed_m3[4] , \speed_m3[5] , \speed_m3[6] , 
            \speed_m3[7] , \speed_m3[8] , \speed_m3[9] , \speed_m3[10] , 
            \speed_m3[11] , \speed_m3[12] , \speed_m3[13] , \speed_m3[14] , 
            \speed_m3[15] , \speed_m3[16] , \speed_m3[17] , \speed_m3[18] , 
            \speed_m3[19] , GND_net, n22097);
    output \speed_m3[0] ;
    input clk_1mhz;
    output [2:0]hallsense_m3;
    input clkout_c_enable_173;
    input H_A_m3_c;
    input H_B_m3_c;
    input H_C_m3_c;
    input rst;
    output \speed_m3[1] ;
    output \speed_m3[2] ;
    output \speed_m3[3] ;
    output \speed_m3[4] ;
    output \speed_m3[5] ;
    output \speed_m3[6] ;
    output \speed_m3[7] ;
    output \speed_m3[8] ;
    output \speed_m3[9] ;
    output \speed_m3[10] ;
    output \speed_m3[11] ;
    output \speed_m3[12] ;
    output \speed_m3[13] ;
    output \speed_m3[14] ;
    output \speed_m3[15] ;
    output \speed_m3[16] ;
    output \speed_m3[17] ;
    output \speed_m3[18] ;
    output \speed_m3[19] ;
    input GND_net;
    input n22097;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire stable_counting;
    wire [19:0]speedt_19__N_1853;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4557;
    wire [19:0]count_19__N_1873;
    
    wire hall3_lat;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_158, hall3_old;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21339, n21304, hall1_lat, hall2_lat, hall1_old, hall2_old, 
        n19429, n19668, n19806, n19666, n11424, n19772, n19676, 
        n19519;
    wire [6:0]n63;
    
    wire n19400, n11422, n4, n12, stable_counting_N_1935, n4_adj_2131, 
        n21340, n14382, n21367, n18112, n18111, n18110, n18109, 
        n18108, n18107, n18106, n18105, n18104, n18103, n18691, 
        n19630, clk_1mhz_enable_179, n19, n24, n20, n22, n16, 
        n21323;
    
    FD1P3AX speed__i1 (.D(speedt_19__N_1853[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_19__N_1873[0]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX speedt_i0_i0 (.D(count_19__N_1873[0]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    LUT4 i2488_2_lut_rep_323_3_lut_4_lut (.A(stable_count[3]), .B(n21339), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21304)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2488_2_lut_rep_323_3_lut_4_lut.init = 16'h78f0;
    FD1P3AX hall1_lat_57 (.D(H_A_m3_c), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m3_c), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m3_c), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(rst), .CK(clk_1mhz), .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(rst), .CK(clk_1mhz), .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n19429), .B(n19668), .C(n19806), .D(n19666), .Z(n11424)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0002;
    LUT4 i16282_2_lut (.A(count[11]), .B(count[14]), .Z(n19668)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16282_2_lut.init = 16'heeee;
    LUT4 i16415_4_lut (.A(count[18]), .B(n19772), .C(n19676), .D(count[16]), 
         .Z(n19806)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16415_4_lut.init = 16'hfffe;
    LUT4 i16280_3_lut (.A(count[12]), .B(count[4]), .C(count[15]), .Z(n19666)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16280_3_lut.init = 16'hfefe;
    LUT4 i16383_4_lut (.A(count[5]), .B(count[7]), .C(count[6]), .D(count[17]), 
         .Z(n19772)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16383_4_lut.init = 16'hfffe;
    LUT4 i16290_2_lut (.A(count[1]), .B(count[19]), .Z(n19676)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16290_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(n19519), .B(stable_count[0]), .C(n63[4]), .D(n19400), 
         .Z(n11422)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_adj_40 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_40.init = 16'h7bde;
    LUT4 i2460_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2460_2_lut.init = 16'h6666;
    LUT4 i6_4_lut (.A(count[10]), .B(n12), .C(count[9]), .D(count[2]), 
         .Z(n19429)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[3]), .B(count[8]), .C(count[13]), .D(count[0]), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i2246_2_lut (.A(stable_counting), .B(stable_counting_N_1935), .Z(n4557)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2246_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_41 (.A(n63[2]), .B(n19519), .C(n63[4]), .D(n4_adj_2131), 
         .Z(stable_counting_N_1935)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_41.init = 16'h0004;
    LUT4 i11814_3_lut (.A(stable_counting), .B(n21340), .C(stable_counting_N_1935), 
         .Z(n14382)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i11814_3_lut.init = 16'ha8a8;
    FD1P3AX speed__i2 (.D(speedt_19__N_1853[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1853[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1853[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1853[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1853[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1853[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1853[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1853[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1853[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1853[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1853[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1853[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1853[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1853[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1853[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1853[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1853[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1853[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1853[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(count_19__N_1873[1]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_1873[2]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_1873[3]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_1873[4]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_1873[5]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_1873[6]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_1873[7]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_1873[8]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_1873[9]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_1873[10]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_1873[11]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_1873[12]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_1873[13]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_1873[14]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_1873[15]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_1873[16]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_1873[17]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_1873[18]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_1873[19]), .CK(clk_1mhz), .CD(n4557), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_1873[1]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[0]), 
         .D(speedt[0]), .Z(speedt_19__N_1853[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[1]), 
         .D(speedt[1]), .Z(speedt_19__N_1853[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX speedt_i0_i2 (.D(count_19__N_1873[2]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_1873[3]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_1873[4]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_1873[5]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_1873[6]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_1873[7]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_1873[8]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_1873[9]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_1873[10]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_1873[11]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_1873[12]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_1873[13]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_1873[14]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_1873[15]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_1873[16]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_1873[17]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_1873[18]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_1873[19]), .SP(clk_1mhz_enable_158), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[2]), 
         .D(speedt[2]), .Z(speedt_19__N_1853[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[3]), 
         .D(speedt[3]), .Z(speedt_19__N_1853[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2481_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21367), .C(stable_count[4]), 
         .D(stable_count[3]), .Z(n63[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2481_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[4]), 
         .D(speedt[4]), .Z(speedt_19__N_1853[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i11515_4_lut (.A(n11424), .B(n11422), .C(stable_counting), .D(stable_counting_N_1935), 
         .Z(clk_1mhz_enable_158)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11515_4_lut.init = 16'hcaea;
    LUT4 i2_3_lut_rep_359 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(n21340)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_359.init = 16'hdede;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[5]), 
         .D(speedt[5]), .Z(speedt_19__N_1853[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[6]), 
         .D(speedt[6]), .Z(speedt_19__N_1853[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .D(n63[1]), 
         .Z(n19519)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[7]), 
         .D(speedt[7]), .Z(speedt_19__N_1853[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[8]), 
         .D(speedt[8]), .Z(speedt_19__N_1853[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[9]), 
         .D(speedt[9]), .Z(speedt_19__N_1853[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[10]), 
         .D(speedt[10]), .Z(speedt_19__N_1853[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[11]), 
         .D(speedt[11]), .Z(speedt_19__N_1853[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[12]), 
         .D(speedt[12]), .Z(speedt_19__N_1853[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[13]), 
         .D(speedt[13]), .Z(speedt_19__N_1853[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[14]), 
         .D(speedt[14]), .Z(speedt_19__N_1853[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[15]), 
         .D(speedt[15]), .Z(speedt_19__N_1853[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[16]), 
         .D(speedt[16]), .Z(speedt_19__N_1853[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[17]), 
         .D(speedt[17]), .Z(speedt_19__N_1853[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[18]), 
         .D(speedt[18]), .Z(speedt_19__N_1853[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11424), .B(n11422), .C(count_19__N_1873[19]), 
         .D(speedt[19]), .Z(speedt_19__N_1853[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18112), 
          .S0(count_19__N_1873[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18111), .COUT(n18112), .S0(count_19__N_1873[17]), .S1(count_19__N_1873[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18110), .COUT(n18111), .S0(count_19__N_1873[15]), .S1(count_19__N_1873[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18109), .COUT(n18110), .S0(count_19__N_1873[13]), .S1(count_19__N_1873[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18108), .COUT(n18109), .S0(count_19__N_1873[11]), .S1(count_19__N_1873[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18107), .COUT(n18108), .S0(count_19__N_1873[9]), .S1(count_19__N_1873[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18106), 
          .COUT(n18107), .S0(count_19__N_1873[7]), .S1(count_19__N_1873[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18105), 
          .COUT(n18106), .S0(count_19__N_1873[5]), .S1(count_19__N_1873[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18104), 
          .COUT(n18105), .S0(count_19__N_1873[3]), .S1(count_19__N_1873[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18103), 
          .COUT(n18104), .S0(count_19__N_1873[1]), .S1(count_19__N_1873[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18103), 
          .S1(count_19__N_1873[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i17197_4_lut (.A(n18691), .B(n19630), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_179)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17197_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_42 (.A(n19), .B(n19429), .C(n24), .D(n20), .Z(n18691)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_42.init = 16'hfffb;
    LUT4 i16245_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19630)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16245_4_lut.init = 16'h7bde;
    LUT4 i6_2_lut (.A(count[17]), .B(count[11]), .Z(n19)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i11_4_lut (.A(count[5]), .B(n22), .C(n16), .D(count[16]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut (.A(count[14]), .B(count[19]), .C(count[6]), .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i9_4_lut (.A(count[18]), .B(count[12]), .C(count[4]), .D(count[7]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[15]), .B(count[1]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i2458_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2458_1_lut.init = 16'h5555;
    LUT4 i2462_2_lut_rep_386 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21367)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2462_2_lut_rep_386.init = 16'h8888;
    LUT4 i2467_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2467_2_lut_3_lut.init = 16'h7878;
    LUT4 i2469_2_lut_rep_358_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21339)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2469_2_lut_rep_358_3_lut.init = 16'h8080;
    LUT4 i2476_2_lut_rep_342_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21323)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2476_2_lut_rep_342_3_lut_4_lut.init = 16'h8000;
    LUT4 i2474_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2474_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21304), .SP(stable_counting), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n63[4]), .SP(stable_counting), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_43 (.A(n63[6]), .B(n63[3]), .C(n21304), .D(n63[2]), 
         .Z(n19400)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_43.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_44 (.A(n63[6]), .B(n63[3]), .C(n21304), .D(stable_count[0]), 
         .Z(n4_adj_2131)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_44.init = 16'hfeff;
    FD1P3IX stable_counting_62 (.D(n22097), .SP(clk_1mhz_enable_179), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14382), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=336, LSE_RLINE=336 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    LUT4 i2495_3_lut_4_lut (.A(stable_count[4]), .B(n21323), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2495_3_lut_4_lut.init = 16'h7f80;
    
endmodule
//
// Verilog Description of module HALL
//

module HALL (clk_1mhz, \speed_m4[0] , hallsense_m4, clkout_c_enable_172, 
            clkout_c_enable_173, HALL_A_OUT_c_c, HALL_B_OUT_c_c, rst, 
            HALL_C_OUT_c_c, \speed_m4[1] , \speed_m4[2] , \speed_m4[3] , 
            \speed_m4[4] , \speed_m4[5] , \speed_m4[6] , \speed_m4[7] , 
            \speed_m4[8] , \speed_m4[9] , \speed_m4[10] , \speed_m4[11] , 
            \speed_m4[12] , \speed_m4[13] , \speed_m4[14] , \speed_m4[15] , 
            \speed_m4[16] , \speed_m4[17] , \speed_m4[18] , \speed_m4[19] , 
            GND_net, n22097);
    input clk_1mhz;
    output \speed_m4[0] ;
    output [2:0]hallsense_m4;
    input clkout_c_enable_172;
    input clkout_c_enable_173;
    input HALL_A_OUT_c_c;
    input HALL_B_OUT_c_c;
    input rst;
    input HALL_C_OUT_c_c;
    output \speed_m4[1] ;
    output \speed_m4[2] ;
    output \speed_m4[3] ;
    output \speed_m4[4] ;
    output \speed_m4[5] ;
    output \speed_m4[6] ;
    output \speed_m4[7] ;
    output \speed_m4[8] ;
    output \speed_m4[9] ;
    output \speed_m4[10] ;
    output \speed_m4[11] ;
    output \speed_m4[12] ;
    output \speed_m4[13] ;
    output \speed_m4[14] ;
    output \speed_m4[15] ;
    output \speed_m4[16] ;
    output \speed_m4[17] ;
    output \speed_m4[18] ;
    output \speed_m4[19] ;
    input GND_net;
    input n22097;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire n18695, n19628, hall3_old, hall3_lat, clk_1mhz_enable_178, 
        n21, n19406, n26, n22, hall1_old, hall2_old, hall1_lat, 
        hall2_lat;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n19658;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21332, n21302, n24, n19614;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_44;
    wire [19:0]count_19__N_1873;
    
    wire n21331, stable_counting, stable_counting_N_1935, n14392, n4565;
    wire [19:0]speedt_19__N_1853;
    
    wire n4;
    wire [6:0]n63;
    
    wire n19522, n11419, n11417, n21350, n21306, n21307, n21349, 
        n18122, n18121, n21319, n18120, n18119, n18118, n18117, 
        n18116, n18115, n18114, n18113, n9, n8, n19798, n19752, 
        n19750, n19403, n21300, n4_adj_2130;
    
    LUT4 i17195_4_lut (.A(n18695), .B(n19628), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_178)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17195_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut (.A(n21), .B(n19406), .C(n26), .D(n22), .Z(n18695)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i16243_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19628)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16243_4_lut.init = 16'h7bde;
    LUT4 i7_4_lut (.A(count[14]), .B(count[8]), .C(n19658), .D(count[9]), 
         .Z(n21)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i2538_2_lut_rep_321_3_lut_4_lut (.A(stable_count[3]), .B(n21332), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21302)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2538_2_lut_rep_321_3_lut_4_lut.init = 16'h78f0;
    LUT4 i12_4_lut (.A(count[1]), .B(n24), .C(n19614), .D(count[11]), 
         .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut.init = 16'hfffe;
    FD1P3AX speedt_i0_i0 (.D(count_19__N_1873[0]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    LUT4 i8_4_lut (.A(count[6]), .B(count[5]), .C(count[18]), .D(count[16]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i16272_2_lut (.A(count[3]), .B(count[13]), .Z(n19658)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16272_2_lut.init = 16'h8888;
    LUT4 i16365_3_lut (.A(n21331), .B(stable_counting), .C(stable_counting_N_1935), 
         .Z(n14392)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16365_3_lut.init = 16'hc8c8;
    FD1S3IX count__i0 (.D(count_19__N_1873[0]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_1853[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_172), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(HALL_A_OUT_c_c), .SP(clkout_c_enable_173), 
            .CK(clk_1mhz), .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    LUT4 i2_3_lut_rep_350 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(n21331)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_350.init = 16'hdede;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4), .C(hall3_lat), .D(n63[1]), 
         .Z(n19522)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    FD1P3AX hall2_lat_58 (.D(HALL_B_OUT_c_c), .SP(clkout_c_enable_173), 
            .CK(clk_1mhz), .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[0]), 
         .D(speedt[0]), .Z(speedt_19__N_1853[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_173), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    LUT4 i2531_2_lut_rep_325_3_lut_4_lut (.A(stable_count[2]), .B(n21350), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21306)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2531_2_lut_rep_325_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2533_2_lut_rep_326_3_lut_4_lut (.A(stable_count[2]), .B(n21350), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21307)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2533_2_lut_rep_326_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[1]), 
         .D(speedt[1]), .Z(speedt_19__N_1853[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[2]), 
         .D(speedt[2]), .Z(speedt_19__N_1853[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[3]), 
         .D(speedt[3]), .Z(speedt_19__N_1853[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX hall3_lat_59 (.D(HALL_C_OUT_c_c), .SP(rst), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(rst), .CK(clk_1mhz), .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[4]), 
         .D(speedt[4]), .Z(speedt_19__N_1853[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[5]), 
         .D(speedt[5]), .Z(speedt_19__N_1853[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[6]), 
         .D(speedt[6]), .Z(speedt_19__N_1853[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[7]), 
         .D(speedt[7]), .Z(speedt_19__N_1853[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX speedt_i0_i19 (.D(count_19__N_1873[19]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[8]), 
         .D(speedt[8]), .Z(speedt_19__N_1853[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[9]), 
         .D(speedt[9]), .Z(speedt_19__N_1853[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX speedt_i0_i18 (.D(count_19__N_1873[18]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_1873[17]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_1873[16]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_1873[15]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_1873[14]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_1873[13]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_1873[12]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_1873[11]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_1873[10]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_1873[9]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_1873[8]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_1873[7]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_1873[6]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_1873[5]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_1873[4]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_1873[3]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_1873[2]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_1873[1]), .SP(clk_1mhz_enable_44), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[10]), 
         .D(speedt[10]), .Z(speedt_19__N_1853[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[11]), 
         .D(speedt[11]), .Z(speedt_19__N_1853[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[12]), 
         .D(speedt[12]), .Z(speedt_19__N_1853[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[13]), 
         .D(speedt[13]), .Z(speedt_19__N_1853[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[14]), 
         .D(speedt[14]), .Z(speedt_19__N_1853[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[15]), 
         .D(speedt[15]), .Z(speedt_19__N_1853[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2251_2_lut (.A(stable_counting), .B(stable_counting_N_1935), .Z(n4565)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2251_2_lut.init = 16'h8888;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[16]), 
         .D(speedt[16]), .Z(speedt_19__N_1853[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[17]), 
         .D(speedt[17]), .Z(speedt_19__N_1853[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[18]), 
         .D(speedt[18]), .Z(speedt_19__N_1853[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX count__i1 (.D(count_19__N_1873[1]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_1873[2]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_1873[3]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_1873[4]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_1873[5]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_1873[6]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_1873[7]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_1873[8]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_1873[9]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_1873[10]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_1873[11]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_1873[12]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_1873[13]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_1873[14]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_1873[15]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_1873[16]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_1873[17]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_1873[18]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_1873[19]), .CK(clk_1mhz), .CD(n4565), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3AX speed__i2 (.D(speedt_19__N_1853[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_1853[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_1853[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_1853[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_1853[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_1853[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_1853[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_1853[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_1853[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_1853[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_1853[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_1853[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_1853[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_1853[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_1853[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_1853[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_1853[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_1853[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_1853[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11419), .B(n11417), .C(count_19__N_1873[19]), 
         .D(speedt[19]), .Z(speedt_19__N_1853[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16227_2_lut_rep_368 (.A(count[4]), .B(count[7]), .Z(n21349)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16227_2_lut_rep_368.init = 16'heeee;
    LUT4 i10_3_lut_4_lut (.A(count[4]), .B(count[7]), .C(count[19]), .D(count[17]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2512_2_lut_rep_369 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21350)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2512_2_lut_rep_369.init = 16'h8888;
    LUT4 i2517_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2517_2_lut_3_lut.init = 16'h7878;
    LUT4 i2524_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2524_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18122), 
          .S0(count_19__N_1873[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18121), .COUT(n18122), .S0(count_19__N_1873[17]), .S1(count_19__N_1873[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    LUT4 i2519_2_lut_rep_351_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21332)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2519_2_lut_rep_351_3_lut.init = 16'h8080;
    LUT4 i2526_2_lut_rep_338_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21319)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2526_2_lut_rep_338_3_lut_4_lut.init = 16'h8000;
    LUT4 i2508_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2508_1_lut.init = 16'h5555;
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18120), .COUT(n18121), .S0(count_19__N_1873[15]), .S1(count_19__N_1873[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18119), .COUT(n18120), .S0(count_19__N_1873[13]), .S1(count_19__N_1873[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18118), .COUT(n18119), .S0(count_19__N_1873[11]), .S1(count_19__N_1873[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18117), .COUT(n18118), .S0(count_19__N_1873[9]), .S1(count_19__N_1873[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    LUT4 i11517_4_lut (.A(n11419), .B(n11417), .C(stable_counting), .D(stable_counting_N_1935), 
         .Z(clk_1mhz_enable_44)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11517_4_lut.init = 16'hcaea;
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18116), 
          .COUT(n18117), .S0(count_19__N_1873[7]), .S1(count_19__N_1873[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18115), 
          .COUT(n18116), .S0(count_19__N_1873[5]), .S1(count_19__N_1873[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18114), 
          .COUT(n18115), .S0(count_19__N_1873[3]), .S1(count_19__N_1873[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18113), 
          .COUT(n18114), .S0(count_19__N_1873[1]), .S1(count_19__N_1873[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18113), 
          .S1(count_19__N_1873[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i5_4_lut (.A(n9), .B(count[9]), .C(n8), .D(count[3]), .Z(n11419)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i3_4_lut (.A(n19406), .B(n21349), .C(n19798), .D(n19752), .Z(n9)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut.init = 16'h0002;
    LUT4 i2_2_lut (.A(count[13]), .B(count[8]), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i16407_4_lut (.A(n19750), .B(count[14]), .C(n19614), .D(count[11]), 
         .Z(n19798)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16407_4_lut.init = 16'hfffe;
    LUT4 i16363_3_lut (.A(count[17]), .B(count[16]), .C(count[1]), .Z(n19752)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16363_3_lut.init = 16'hfefe;
    LUT4 i16361_4_lut (.A(count[18]), .B(count[6]), .C(count[5]), .D(count[19]), 
         .Z(n19750)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16361_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n19522), .B(stable_count[0]), .C(n21306), .D(n19403), 
         .Z(n11417)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_adj_37 (.A(n63[2]), .B(n19522), .C(n21300), .D(n4_adj_2130), 
         .Z(stable_counting_N_1935)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_37.init = 16'h0004;
    FD1P3IX stable_counting_62 (.D(n22097), .SP(clk_1mhz_enable_178), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21302), .SP(stable_counting), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21306), .SP(stable_counting), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_38 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_38.init = 16'h7bde;
    LUT4 i2510_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2510_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_4_lut_adj_39 (.A(n63[3]), .B(n63[6]), .C(n21302), .D(n63[2]), 
         .Z(n19403)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_2_lut_4_lut_adj_39.init = 16'hfffe;
    LUT4 i16229_2_lut (.A(count[12]), .B(count[15]), .Z(n19614)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16229_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(count[10]), .B(count[2]), .C(count[0]), .Z(n19406)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14392), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=346, LSE_RLINE=346 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_319_4_lut (.A(stable_count[5]), .B(n21307), .C(n63[6]), 
         .D(n63[3]), .Z(n21300)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_319_4_lut.init = 16'hfff6;
    LUT4 i2545_3_lut_4_lut (.A(stable_count[4]), .B(n21319), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2545_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21332), .C(stable_count[0]), 
         .D(stable_count[4]), .Z(n4_adj_2130)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h7f8f;
    
endmodule
