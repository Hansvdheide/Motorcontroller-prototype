// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.8.0.115.3
// Netlist written on Fri Jun 30 13:54:24 2017
//
// Verilog Description of module SPI_loopback_Top
//

module SPI_loopback_Top (CS, SCK, MOSI, MISO, HALL_A_OUT, HALL_B_OUT, 
            HALL_C_OUT, LED1, LED2, LED3, LED4, clkout, H_A_m1, 
            H_B_m1, H_C_m1, MA_m1, MB_m1, MC_m1, H_A_m2, H_B_m2, 
            H_C_m2, MA_m2, MB_m2, MC_m2, H_A_m3, H_B_m3, H_C_m3, 
            MA_m3, MB_m3, MC_m3, H_A_m4, H_B_m4, H_C_m4, MA_m4, 
            MB_m4, MC_m4);   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(24[8:24])
    input CS;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(27[2:4])
    input SCK;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(28[2:5])
    input MOSI;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(29[2:6])
    output MISO;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(30[2:6])
    output HALL_A_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(33[2:12])
    output HALL_B_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(34[2:12])
    output HALL_C_OUT;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(35[2:12])
    output LED1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(38[2:6])
    output LED2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(39[2:6])
    output LED3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(40[2:6])
    output LED4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(41[2:6])
    output clkout;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    input H_A_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(47[2:8])
    input H_B_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(48[2:8])
    input H_C_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(49[2:8])
    output [1:0]MA_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    output [1:0]MB_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    output [1:0]MC_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    input H_A_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(55[2:8])
    input H_B_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(56[2:8])
    input H_C_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(57[2:8])
    output [1:0]MA_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    output [1:0]MB_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    output [1:0]MC_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    input H_A_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(63[2:8])
    input H_B_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(64[2:8])
    input H_C_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(65[2:8])
    output [1:0]MA_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    output [1:0]MB_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    output [1:0]MC_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    input H_A_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(71[2:8])
    input H_B_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(72[2:8])
    input H_C_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(73[2:8])
    output [1:0]MA_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    output [1:0]MB_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    output [1:0]MC_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    wire clk_N_875 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    
    wire GND_net, VCC_net, CS_c, SCK_c, MOSI_c, HALL_A_OUT_c_c, 
        HALL_B_OUT_c_c, HALL_C_OUT_c_c, LED1_c, LED2_c, LED3_c, LED4_c, 
        MA_m1_c_1, MA_m1_c_0, MB_m1_c_1, MB_m1_c_0, MC_m1_c_1, MC_m1_c_0, 
        H_A_m2_c, H_B_m2_c, H_C_m2_c, MA_m2_c_1, MA_m2_c_0, MB_m2_c_1, 
        MB_m2_c_0, MC_m2_c_1, MC_m2_c_0, H_A_m3_c, H_B_m3_c, H_C_m3_c, 
        MA_m3_c_1, MA_m3_c_0, MB_m3_c_1, MB_m3_c_0, MC_m3_c_1, MC_m3_c_0, 
        H_A_m4_c, H_B_m4_c, H_C_m4_c, MA_m4_c_1, MA_m4_c_0, MB_m4_c_1, 
        MB_m4_c_0, MC_m4_c_1, MC_m4_c_0, rst, enable_m1, enable_m2, 
        enable_m3, enable_m4;
    wire [20:0]speed_set_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(99[9:21])
    wire [20:0]speed_set_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(100[9:21])
    wire [20:0]speed_set_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(101[9:21])
    wire [20:0]speed_set_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(102[9:21])
    wire [20:0]speed_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(104[9:17])
    wire [20:0]speed_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(105[9:17])
    wire [20:0]speed_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(106[9:17])
    wire [20:0]speed_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(107[9:17])
    wire [2:0]hallsense_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(110[9:21])
    wire [2:0]hallsense_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(111[9:21])
    wire [2:0]hallsense_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(112[9:21])
    wire [2:0]hallsense_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(113[9:21])
    
    wire PWM_m1, PWM_m2, PWM_m3, PWM_m4;
    wire [9:0]PWMdut_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(120[9:18])
    wire [9:0]PWMdut_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(121[9:18])
    wire [9:0]PWMdut_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(122[9:18])
    wire [9:0]PWMdut_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(123[9:18])
    
    wire dir_m1, dir_m2, dir_m3, dir_m4;
    wire [13:0]start_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(135[9:18])
    wire [20:0]speed_avg_m1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(144[9:21])
    wire [20:0]speed_avg_m2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(145[9:21])
    wire [20:0]speed_avg_m3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(146[9:21])
    wire [20:0]speed_avg_m4;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(147[9:21])
    
    wire n18657, n4530, n4531, n3241, n3207, n3139, n3105, n3037, 
        n3003, n2935, MISO_N_816, n4520, n4504, n4497, n4494, 
        n4492, n4491, n2901, n4510, n4511, n4512, n21422, n4513, 
        n4514, n4515, n4516, n4517, n4519, n4522;
    wire [25:0]subOut_24__N_1369;
    
    wire n14195, n4527, n4528, n4529, n4525, n4499, n4489, n4488, 
        n4487, n4521, n4518, n4503, n4486, n4485, n4500, n4501, 
        n4502, n4505, n4506, n4526, n4523, n4524, n18370, n18369, 
        n18368, n18367, n18366, n18365, n18364, n6, n4493, n4495, 
        n4496, n4498, n4490, n4484, n19649, n62, n63, n64, n65, 
        n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
        n5199, n10485, n18732, n18749, n14203, clkout_c_enable_360, 
        clkout_c_enable_362, clkout_c_enable_266, n22211, n22206, n14208, 
        n21487, n21485, n21484, n21476, n14200, n21453, n21452, 
        n21451, n21449;
    
    VHI i2 (.Z(VCC_net));
    OSCH OSCInst0 (.STDBY(GND_net), .OSC(clkout_c)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCInst0.NOM_FREQ = "38.00";
    FD1S3AX rst_12 (.D(n21422), .CK(clkout_c), .Q(rst));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(386[3] 393[10])
    defparam rst_12.GSR = "DISABLED";
    GSR GSR_INST (.GSR(n22211));
    LUT4 m1_lut (.Z(n22206)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    OB MA_m2_pad_0 (.I(MA_m2_c_0), .O(MA_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    FD1P3AX start_cnt_2121__i0 (.D(n75), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i0.GSR = "DISABLED";
    OB HALL_B_OUT_pad (.I(HALL_B_OUT_c_c), .O(HALL_B_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(34[2:12])
    OB HALL_A_OUT_pad (.I(HALL_A_OUT_c_c), .O(HALL_A_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(33[2:12])
    OB MA_m2_pad_1 (.I(MA_m2_c_1), .O(MA_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(58[2:7])
    IB HALL_B_OUT_c_pad (.I(H_B_m1), .O(HALL_B_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(48[2:8])
    OBZ n5198_pad (.I(MISO_N_816), .T(n5199), .O(MISO));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    IB HALL_A_OUT_c_pad (.I(H_A_m1), .O(HALL_A_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(47[2:8])
    IB MOSI_pad (.I(MOSI), .O(MOSI_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(29[2:6])
    IB SCK_pad (.I(SCK), .O(SCK_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(28[2:5])
    IB CS_pad (.I(CS), .O(CS_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(27[2:4])
    OB MC_m4_pad_0 (.I(MC_m4_c_0), .O(MC_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    OB MC_m4_pad_1 (.I(MC_m4_c_1), .O(MC_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(76[2:7])
    OB MB_m4_pad_0 (.I(MB_m4_c_0), .O(MB_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    OB MB_m4_pad_1 (.I(MB_m4_c_1), .O(MB_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(75[2:7])
    OB MC_m1_pad_0 (.I(MC_m1_c_0), .O(MC_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    OB MC_m1_pad_1 (.I(MC_m1_c_1), .O(MC_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(52[2:7])
    OB MA_m4_pad_0 (.I(MA_m4_c_0), .O(MA_m4[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_0 (.I(MB_m1_c_0), .O(MB_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    OB MA_m4_pad_1 (.I(MA_m4_c_1), .O(MA_m4[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(74[2:7])
    OB MB_m1_pad_1 (.I(MB_m1_c_1), .O(MB_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(51[2:7])
    OB MC_m3_pad_0 (.I(MC_m3_c_0), .O(MC_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    IB H_C_m4_pad (.I(H_C_m4), .O(H_C_m4_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(73[2:8])
    OB MA_m1_pad_0 (.I(MA_m1_c_0), .O(MA_m1[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    OB MC_m3_pad_1 (.I(MC_m3_c_1), .O(MC_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(68[2:7])
    IB H_B_m4_pad (.I(H_B_m4), .O(H_B_m4_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(72[2:8])
    LUT4 mux_2193_i1_3_lut (.A(n4506), .B(n4531), .C(n19649), .Z(subOut_24__N_1369[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i1_3_lut.init = 16'hacac;
    OB MA_m1_pad_1 (.I(MA_m1_c_1), .O(MA_m1[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(50[2:7])
    OB MB_m3_pad_0 (.I(MB_m3_c_0), .O(MB_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    IB H_A_m4_pad (.I(H_A_m4), .O(H_A_m4_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(71[2:8])
    OB clkout_pad (.I(clkout_c), .O(clkout));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    OB MB_m3_pad_1 (.I(MB_m3_c_1), .O(MB_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(67[2:7])
    IB H_C_m3_pad (.I(H_C_m3), .O(H_C_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(65[2:8])
    OB LED4_pad (.I(LED4_c), .O(LED4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(41[2:6])
    OB MA_m3_pad_0 (.I(MA_m3_c_0), .O(MA_m3[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    IB H_B_m3_pad (.I(H_B_m3), .O(H_B_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(64[2:8])
    OB LED3_pad (.I(LED3_c), .O(LED3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(40[2:6])
    OB MA_m3_pad_1 (.I(MA_m3_c_1), .O(MA_m3[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(66[2:7])
    IB H_A_m3_pad (.I(H_A_m3), .O(H_A_m3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(63[2:8])
    OB LED2_pad (.I(LED2_c), .O(LED2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(39[2:6])
    OB MC_m2_pad_0 (.I(MC_m2_c_0), .O(MC_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    IB H_C_m2_pad (.I(H_C_m2), .O(H_C_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(57[2:8])
    OB LED1_pad (.I(LED1_c), .O(LED1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(38[2:6])
    OB MC_m2_pad_1 (.I(MC_m2_c_1), .O(MC_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(60[2:7])
    IB H_B_m2_pad (.I(H_B_m2), .O(H_B_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(56[2:8])
    OB HALL_C_OUT_pad (.I(HALL_C_OUT_c_c), .O(HALL_C_OUT));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(35[2:12])
    OB MB_m2_pad_0 (.I(MB_m2_c_0), .O(MB_m2[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    IB H_A_m2_pad (.I(H_A_m2), .O(H_A_m2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(55[2:8])
    OB MB_m2_pad_1 (.I(MB_m2_c_1), .O(MB_m2[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(59[2:7])
    IB HALL_C_OUT_c_pad (.I(H_C_m1), .O(HALL_C_OUT_c_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(49[2:8])
    LUT4 i8004_4_lut_rep_348 (.A(n21484), .B(hallsense_m4[2]), .C(dir_m4), 
         .D(hallsense_m4[0]), .Z(n21449)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i8004_4_lut_rep_348.init = 16'h755d;
    LUT4 i11602_1_lut_4_lut (.A(n21484), .B(hallsense_m4[2]), .C(dir_m4), 
         .D(hallsense_m4[0]), .Z(n14208)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i11602_1_lut_4_lut.init = 16'h8aa2;
    LUT4 i7993_4_lut_rep_350 (.A(n21476), .B(hallsense_m1[2]), .C(dir_m1), 
         .D(hallsense_m1[0]), .Z(n21451)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i7993_4_lut_rep_350.init = 16'h755d;
    LUT4 i11589_1_lut_4_lut (.A(n21476), .B(hallsense_m1[2]), .C(dir_m1), 
         .D(hallsense_m1[0]), .Z(n14195)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i11589_1_lut_4_lut.init = 16'h8aa2;
    LUT4 i8001_4_lut_rep_351 (.A(n21485), .B(hallsense_m3[2]), .C(dir_m3), 
         .D(hallsense_m3[0]), .Z(n21452)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i8001_4_lut_rep_351.init = 16'h755d;
    LUT4 i11597_1_lut_4_lut (.A(n21485), .B(hallsense_m3[2]), .C(dir_m3), 
         .D(hallsense_m3[0]), .Z(n14203)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i11597_1_lut_4_lut.init = 16'h8aa2;
    LUT4 i7998_4_lut_rep_352 (.A(n21487), .B(hallsense_m2[2]), .C(dir_m2), 
         .D(hallsense_m2[0]), .Z(n21453)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i7998_4_lut_rep_352.init = 16'h755d;
    LUT4 i11594_1_lut_4_lut (.A(n21487), .B(hallsense_m2[2]), .C(dir_m2), 
         .D(hallsense_m2[0]), .Z(n14200)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i11594_1_lut_4_lut.init = 16'h8aa2;
    LUT4 i3_4_lut (.A(n18732), .B(start_cnt[10]), .C(start_cnt[9]), .D(start_cnt[8]), 
         .Z(n18657)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_191 (.A(n18749), .B(n6), .C(start_cnt[6]), .D(start_cnt[4]), 
         .Z(n18732)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_191.init = 16'hfefc;
    LUT4 i3_4_lut_adj_192 (.A(start_cnt[0]), .B(start_cnt[3]), .C(start_cnt[2]), 
         .D(start_cnt[1]), .Z(n18749)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_192.init = 16'hfffe;
    LUT4 i2_2_lut (.A(start_cnt[7]), .B(start_cnt[5]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 mux_2193_i18_3_lut (.A(n4489), .B(n4514), .C(n19649), .Z(subOut_24__N_1369[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i18_3_lut.init = 16'hacac;
    LUT4 mux_2193_i19_3_lut (.A(n4488), .B(n4513), .C(n19649), .Z(subOut_24__N_1369[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i19_3_lut.init = 16'hacac;
    LUT4 mux_2193_i20_3_lut (.A(n4487), .B(n4512), .C(n19649), .Z(subOut_24__N_1369[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i20_3_lut.init = 16'hacac;
    LUT4 mux_2193_i21_3_lut (.A(n4486), .B(n4511), .C(n19649), .Z(subOut_24__N_1369[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i21_3_lut.init = 16'hacac;
    LUT4 mux_2193_i22_3_lut (.A(n4485), .B(n4510), .C(n19649), .Z(subOut_24__N_1369[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i22_3_lut.init = 16'hacac;
    LUT4 mux_2193_i25_3_lut (.A(n4484), .B(n4510), .C(n19649), .Z(subOut_24__N_1369[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i25_3_lut.init = 16'hacac;
    LUT4 i2388_4_lut_rep_321 (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18657), .Z(n21422)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2388_4_lut_rep_321.init = 16'hccc8;
    LUT4 i9378_1_lut_4_lut (.A(start_cnt[12]), .B(start_cnt[13]), .C(start_cnt[11]), 
         .D(n18657), .Z(clkout_c_enable_360)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i9378_1_lut_4_lut.init = 16'h3337;
    LUT4 i7981_2_lut (.A(n21422), .B(n62), .Z(n10485)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam i7981_2_lut.init = 16'heeee;
    LUT4 mux_2193_i2_3_lut (.A(n4505), .B(n4530), .C(n19649), .Z(subOut_24__N_1369[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i2_3_lut.init = 16'hacac;
    LUT4 i17220_4_lut (.A(n21484), .B(hallsense_m4[1]), .C(dir_m4), .D(hallsense_m4[0]), 
         .Z(n3241)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i17220_4_lut.init = 16'h8aa2;
    LUT4 i17218_4_lut (.A(n21484), .B(hallsense_m4[2]), .C(dir_m4), .D(hallsense_m4[1]), 
         .Z(n3207)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(128[9:15])
    defparam i17218_4_lut.init = 16'h8aa2;
    LUT4 i17216_4_lut (.A(n21485), .B(hallsense_m3[1]), .C(dir_m3), .D(hallsense_m3[0]), 
         .Z(n3139)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i17216_4_lut.init = 16'h8aa2;
    LUT4 i17214_4_lut (.A(n21485), .B(hallsense_m3[2]), .C(dir_m3), .D(hallsense_m3[1]), 
         .Z(n3105)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(127[9:15])
    defparam i17214_4_lut.init = 16'h8aa2;
    LUT4 i17212_4_lut (.A(n21487), .B(hallsense_m2[1]), .C(dir_m2), .D(hallsense_m2[0]), 
         .Z(n3037)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i17212_4_lut.init = 16'h8aa2;
    LUT4 i17210_4_lut (.A(n21487), .B(hallsense_m2[2]), .C(dir_m2), .D(hallsense_m2[1]), 
         .Z(n3003)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(126[9:15])
    defparam i17210_4_lut.init = 16'h8aa2;
    LUT4 i17208_4_lut (.A(n21476), .B(hallsense_m1[1]), .C(dir_m1), .D(hallsense_m1[0]), 
         .Z(n2935)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i17208_4_lut.init = 16'h8aa2;
    LUT4 i17206_4_lut (.A(n21476), .B(hallsense_m1[2]), .C(dir_m1), .D(hallsense_m1[1]), 
         .Z(n2901)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(125[9:15])
    defparam i17206_4_lut.init = 16'h8aa2;
    CCU2D start_cnt_2121_add_4_15 (.A0(start_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18370), .S0(n62));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_15.INIT0 = 16'hfaaa;
    defparam start_cnt_2121_add_4_15.INIT1 = 16'h0000;
    defparam start_cnt_2121_add_4_15.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_15.INJECT1_1 = "NO";
    CCU2D start_cnt_2121_add_4_13 (.A0(start_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18369), .COUT(n18370), .S0(n64), .S1(n63));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_13.INIT0 = 16'hfaaa;
    defparam start_cnt_2121_add_4_13.INIT1 = 16'hfaaa;
    defparam start_cnt_2121_add_4_13.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_13.INJECT1_1 = "NO";
    CCU2D start_cnt_2121_add_4_11 (.A0(start_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18368), .COUT(n18369), .S0(n66), .S1(n65));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_11.INIT0 = 16'hfaaa;
    defparam start_cnt_2121_add_4_11.INIT1 = 16'hfaaa;
    defparam start_cnt_2121_add_4_11.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_11.INJECT1_1 = "NO";
    CCU2D start_cnt_2121_add_4_9 (.A0(start_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18367), .COUT(n18368), .S0(n68), .S1(n67));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_9.INIT0 = 16'hfaaa;
    defparam start_cnt_2121_add_4_9.INIT1 = 16'hfaaa;
    defparam start_cnt_2121_add_4_9.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_9.INJECT1_1 = "NO";
    CCU2D start_cnt_2121_add_4_7 (.A0(start_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18366), .COUT(n18367), .S0(n70), .S1(n69));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_7.INIT0 = 16'hfaaa;
    defparam start_cnt_2121_add_4_7.INIT1 = 16'hfaaa;
    defparam start_cnt_2121_add_4_7.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_7.INJECT1_1 = "NO";
    CLKDIV CLKDIV_I (.clk_N_875(clk_N_875), .clkout_c(clkout_c), .clk_1mhz(clk_1mhz), 
           .pwm_clk(pwm_clk), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(308[14:20])
    CCU2D start_cnt_2121_add_4_5 (.A0(start_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18365), .COUT(n18366), .S0(n72), .S1(n71));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_5.INIT0 = 16'hfaaa;
    defparam start_cnt_2121_add_4_5.INIT1 = 16'hfaaa;
    defparam start_cnt_2121_add_4_5.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_5.INJECT1_1 = "NO";
    HALL_U4 HALL_I_M2 (.clk_1mhz(clk_1mhz), .\speed_m2[0] (speed_m2[0]), 
            .hallsense_m2({hallsense_m2}), .rst(rst), .H_B_m2_c(H_B_m2_c), 
            .clkout_c_enable_266(clkout_c_enable_266), .H_A_m2_c(H_A_m2_c), 
            .clkout_c_enable_362(clkout_c_enable_362), .H_C_m2_c(H_C_m2_c), 
            .\speed_m2[1] (speed_m2[1]), .\speed_m2[2] (speed_m2[2]), .\speed_m2[3] (speed_m2[3]), 
            .\speed_m2[4] (speed_m2[4]), .\speed_m2[5] (speed_m2[5]), .\speed_m2[6] (speed_m2[6]), 
            .\speed_m2[7] (speed_m2[7]), .\speed_m2[8] (speed_m2[8]), .\speed_m2[9] (speed_m2[9]), 
            .\speed_m2[10] (speed_m2[10]), .\speed_m2[11] (speed_m2[11]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_m2[13] (speed_m2[13]), 
            .\speed_m2[14] (speed_m2[14]), .\speed_m2[15] (speed_m2[15]), 
            .\speed_m2[16] (speed_m2[16]), .\speed_m2[17] (speed_m2[17]), 
            .\speed_m2[18] (speed_m2[18]), .\speed_m2[19] (speed_m2[19]), 
            .GND_net(GND_net), .n22206(n22206));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(332[14:18])
    LUT4 mux_2193_i3_3_lut (.A(n4504), .B(n4529), .C(n19649), .Z(subOut_24__N_1369[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i3_3_lut.init = 16'hacac;
    CCU2D start_cnt_2121_add_4_3 (.A0(start_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18364), .COUT(n18365), .S0(n74), .S1(n73));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_3.INIT0 = 16'hfaaa;
    defparam start_cnt_2121_add_4_3.INIT1 = 16'hfaaa;
    defparam start_cnt_2121_add_4_3.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_3.INJECT1_1 = "NO";
    CCU2D start_cnt_2121_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18364), .S1(n75));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121_add_4_1.INIT0 = 16'hF000;
    defparam start_cnt_2121_add_4_1.INIT1 = 16'h0555;
    defparam start_cnt_2121_add_4_1.INJECT1_0 = "NO";
    defparam start_cnt_2121_add_4_1.INJECT1_1 = "NO";
    LUT4 mux_2193_i4_3_lut (.A(n4503), .B(n4528), .C(n19649), .Z(subOut_24__N_1369[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i4_3_lut.init = 16'hacac;
    COMMUTATION_U7 COM_I_M2 (.MB_m2_c_0(MB_m2_c_0), .clkout_c(clkout_c), 
            .MC_m2_c_0(MC_m2_c_0), .n21487(n21487), .dir_m2(dir_m2), .hallsense_m2({hallsense_m2}), 
            .MA_m2_c_1(MA_m2_c_1), .n21453(n21453), .PWM_m2(PWM_m2), .MC_m2_c_1(MC_m2_c_1), 
            .n3037(n3037), .MB_m2_c_1(MB_m2_c_1), .n3003(n3003), .LED2_c(LED2_c), 
            .enable_m2(enable_m2), .MA_m2_c_0(MA_m2_c_0), .n14200(n14200));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(335[13:24])
    LUT4 mux_2193_i5_3_lut (.A(n4502), .B(n4527), .C(n19649), .Z(subOut_24__N_1369[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i5_3_lut.init = 16'hacac;
    COMMUTATION_U8 COM_I_M1 (.n21476(n21476), .dir_m1(dir_m1), .hallsense_m1({hallsense_m1}), 
            .MA_m1_c_0(MA_m1_c_0), .clkout_c(clkout_c), .n14195(n14195), 
            .MB_m1_c_0(MB_m1_c_0), .MC_m1_c_0(MC_m1_c_0), .MA_m1_c_1(MA_m1_c_1), 
            .n21451(n21451), .LED1_c(LED1_c), .enable_m1(enable_m1), .PWM_m1(PWM_m1), 
            .MC_m1_c_1(MC_m1_c_1), .n2935(n2935), .MB_m1_c_1(MB_m1_c_1), 
            .n2901(n2901));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(325[13:24])
    LUT4 mux_2193_i6_3_lut (.A(n4501), .B(n4526), .C(n19649), .Z(subOut_24__N_1369[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i6_3_lut.init = 16'hacac;
    LUT4 mux_2193_i7_3_lut (.A(n4500), .B(n4525), .C(n19649), .Z(subOut_24__N_1369[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i7_3_lut.init = 16'hacac;
    LUT4 mux_2193_i8_3_lut (.A(n4499), .B(n4524), .C(n19649), .Z(subOut_24__N_1369[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i8_3_lut.init = 16'hacac;
    LUT4 mux_2193_i9_3_lut (.A(n4498), .B(n4523), .C(n19649), .Z(subOut_24__N_1369[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i9_3_lut.init = 16'hacac;
    LUT4 mux_2193_i10_3_lut (.A(n4497), .B(n4522), .C(n19649), .Z(subOut_24__N_1369[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i10_3_lut.init = 16'hacac;
    LUT4 mux_2193_i11_3_lut (.A(n4496), .B(n4521), .C(n19649), .Z(subOut_24__N_1369[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i11_3_lut.init = 16'hacac;
    HALL_U5 HALL_I_M1 (.clk_1mhz(clk_1mhz), .GND_net(GND_net), .\speed_m1[0] (speed_m1[0]), 
            .hallsense_m1({hallsense_m1}), .clkout_c_enable_362(clkout_c_enable_362), 
            .clkout_c_enable_266(clkout_c_enable_266), .HALL_A_OUT_c_c(HALL_A_OUT_c_c), 
            .HALL_B_OUT_c_c(HALL_B_OUT_c_c), .HALL_C_OUT_c_c(HALL_C_OUT_c_c), 
            .\speed_m1[1] (speed_m1[1]), .\speed_m1[2] (speed_m1[2]), .\speed_m1[3] (speed_m1[3]), 
            .\speed_m1[4] (speed_m1[4]), .\speed_m1[5] (speed_m1[5]), .\speed_m1[6] (speed_m1[6]), 
            .\speed_m1[7] (speed_m1[7]), .\speed_m1[8] (speed_m1[8]), .\speed_m1[9] (speed_m1[9]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_m1[11] (speed_m1[11]), 
            .\speed_m1[12] (speed_m1[12]), .\speed_m1[13] (speed_m1[13]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_m1[15] (speed_m1[15]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_m1[17] (speed_m1[17]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_m1[19] (speed_m1[19]), 
            .n22206(n22206));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(322[14:18])
    COMMUTATION_U6 COM_I_M3 (.MB_m3_c_0(MB_m3_c_0), .clkout_c(clkout_c), 
            .MC_m3_c_0(MC_m3_c_0), .n21485(n21485), .dir_m3(dir_m3), .hallsense_m3({hallsense_m3}), 
            .LED3_c(LED3_c), .enable_m3(enable_m3), .PWM_m3(PWM_m3), .MA_m3_c_1(MA_m3_c_1), 
            .n21452(n21452), .MA_m3_c_0(MA_m3_c_0), .n14203(n14203), .MC_m3_c_1(MC_m3_c_1), 
            .n3139(n3139), .MB_m3_c_1(MB_m3_c_1), .n3105(n3105));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(345[13:24])
    HALL_U3 HALL_I_M3 (.clk_1mhz(clk_1mhz), .\speed_m3[0] (speed_m3[0]), 
            .hallsense_m3({hallsense_m3}), .clkout_c_enable_362(clkout_c_enable_362), 
            .H_A_m3_c(H_A_m3_c), .H_B_m3_c(H_B_m3_c), .H_C_m3_c(H_C_m3_c), 
            .\speed_m3[1] (speed_m3[1]), .\speed_m3[2] (speed_m3[2]), .\speed_m3[3] (speed_m3[3]), 
            .\speed_m3[4] (speed_m3[4]), .\speed_m3[5] (speed_m3[5]), .\speed_m3[6] (speed_m3[6]), 
            .\speed_m3[7] (speed_m3[7]), .\speed_m3[8] (speed_m3[8]), .\speed_m3[9] (speed_m3[9]), 
            .\speed_m3[10] (speed_m3[10]), .\speed_m3[11] (speed_m3[11]), 
            .\speed_m3[12] (speed_m3[12]), .\speed_m3[13] (speed_m3[13]), 
            .\speed_m3[14] (speed_m3[14]), .\speed_m3[15] (speed_m3[15]), 
            .\speed_m3[16] (speed_m3[16]), .\speed_m3[17] (speed_m3[17]), 
            .\speed_m3[18] (speed_m3[18]), .\speed_m3[19] (speed_m3[19]), 
            .GND_net(GND_net), .n22206(n22206));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(342[14:18])
    LUT4 mux_2193_i12_3_lut (.A(n4495), .B(n4520), .C(n19649), .Z(subOut_24__N_1369[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i12_3_lut.init = 16'hacac;
    LUT4 mux_2193_i13_3_lut (.A(n4494), .B(n4519), .C(n19649), .Z(subOut_24__N_1369[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i13_3_lut.init = 16'hacac;
    COMMUTATION COM_I_M4 (.MB_m4_c_0(MB_m4_c_0), .clkout_c(clkout_c), .MC_m4_c_0(MC_m4_c_0), 
            .n21484(n21484), .dir_m4(dir_m4), .hallsense_m4({hallsense_m4}), 
            .PWM_m4(PWM_m4), .MA_m4_c_1(MA_m4_c_1), .n21449(n21449), .LED4_c(LED4_c), 
            .enable_m4(enable_m4), .MC_m4_c_1(MC_m4_c_1), .n3241(n3241), 
            .MB_m4_c_1(MB_m4_c_1), .n3207(n3207), .MA_m4_c_0(MA_m4_c_0), 
            .n14208(n14208));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(355[13:24])
    LUT4 mux_2193_i14_3_lut (.A(n4493), .B(n4518), .C(n19649), .Z(subOut_24__N_1369[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i14_3_lut.init = 16'hacac;
    LUT4 mux_2193_i15_3_lut (.A(n4492), .B(n4517), .C(n19649), .Z(subOut_24__N_1369[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i15_3_lut.init = 16'hacac;
    LUT4 mux_2193_i16_3_lut (.A(n4491), .B(n4516), .C(n19649), .Z(subOut_24__N_1369[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i16_3_lut.init = 16'hacac;
    LUT4 mux_2193_i17_3_lut (.A(n4490), .B(n4515), .C(n19649), .Z(subOut_24__N_1369[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam mux_2193_i17_3_lut.init = 16'hacac;
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    FD1S3AX rst_12_rep_407 (.D(n21422), .CK(clkout_c), .Q(clkout_c_enable_362));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(386[3] 393[10])
    defparam rst_12_rep_407.GSR = "DISABLED";
    AVG_SPEED AVG_SPEED_M4 (.\speed_avg_m4[0] (speed_avg_m4[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m4[0] (speed_m4[0]), .\speed_avg_m4[1] (speed_avg_m4[1]), 
            .\speed_m4[1] (speed_m4[1]), .\speed_avg_m4[2] (speed_avg_m4[2]), 
            .\speed_m4[2] (speed_m4[2]), .\speed_avg_m4[3] (speed_avg_m4[3]), 
            .\speed_m4[3] (speed_m4[3]), .\speed_avg_m4[4] (speed_avg_m4[4]), 
            .\speed_m4[4] (speed_m4[4]), .\speed_avg_m4[5] (speed_avg_m4[5]), 
            .\speed_m4[5] (speed_m4[5]), .\speed_avg_m4[6] (speed_avg_m4[6]), 
            .\speed_m4[6] (speed_m4[6]), .\speed_avg_m4[7] (speed_avg_m4[7]), 
            .\speed_m4[7] (speed_m4[7]), .\speed_avg_m4[8] (speed_avg_m4[8]), 
            .\speed_m4[8] (speed_m4[8]), .\speed_avg_m4[9] (speed_avg_m4[9]), 
            .\speed_m4[9] (speed_m4[9]), .\speed_avg_m4[10] (speed_avg_m4[10]), 
            .\speed_m4[10] (speed_m4[10]), .\speed_avg_m4[11] (speed_avg_m4[11]), 
            .\speed_m4[11] (speed_m4[11]), .\speed_avg_m4[12] (speed_avg_m4[12]), 
            .\speed_m4[12] (speed_m4[12]), .\speed_avg_m4[13] (speed_avg_m4[13]), 
            .\speed_m4[13] (speed_m4[13]), .\speed_avg_m4[14] (speed_avg_m4[14]), 
            .\speed_m4[14] (speed_m4[14]), .\speed_avg_m4[15] (speed_avg_m4[15]), 
            .\speed_m4[15] (speed_m4[15]), .\speed_avg_m4[16] (speed_avg_m4[16]), 
            .\speed_m4[16] (speed_m4[16]), .\speed_avg_m4[17] (speed_avg_m4[17]), 
            .\speed_m4[17] (speed_m4[17]), .\speed_avg_m4[18] (speed_avg_m4[18]), 
            .\speed_m4[18] (speed_m4[18]), .\speed_avg_m4[19] (speed_avg_m4[19]), 
            .\speed_m4[19] (speed_m4[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(370[17:26])
    FD1P3AX start_cnt_2121__i1 (.D(n74), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i1.GSR = "DISABLED";
    FD1S3AX rst_12_rep_406 (.D(n21422), .CK(clkout_c), .Q(clkout_c_enable_266));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(386[3] 393[10])
    defparam rst_12_rep_406.GSR = "DISABLED";
    FD1S3AX rst_12_rep_405 (.D(n21422), .CK(clkout_c), .Q(n22211));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(386[3] 393[10])
    defparam rst_12_rep_405.GSR = "DISABLED";
    SPI SPI_I (.GND_net(GND_net), .clkout_c(clkout_c), .MISO_N_816(MISO_N_816), 
        .n22211(n22211), .speed_set_m2({speed_set_m2}), .speed_set_m4({speed_set_m4}), 
        .speed_set_m1({speed_set_m1}), .enable_m1(enable_m1), .enable_m2(enable_m2), 
        .enable_m3(enable_m3), .enable_m4(enable_m4), .clkout_c_enable_362(clkout_c_enable_362), 
        .CS_c(CS_c), .SCK_c(SCK_c), .MOSI_c(MOSI_c), .clkout_c_enable_266(clkout_c_enable_266), 
        .rst(rst), .n5199(n5199), .speed_set_m3({speed_set_m3}));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(313[10:13])
    FD1P3AX start_cnt_2121__i2 (.D(n73), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i2.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i3 (.D(n72), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i3.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i4 (.D(n71), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i4.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i5 (.D(n70), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i5.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i6 (.D(n69), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i6.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i7 (.D(n68), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i7.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i8 (.D(n67), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i8.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i9 (.D(n66), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i9.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i10 (.D(n65), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i10.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i11 (.D(n64), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i11.GSR = "DISABLED";
    FD1P3AX start_cnt_2121__i12 (.D(n63), .SP(clkout_c_enable_360), .CK(clkout_c), 
            .Q(start_cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i12.GSR = "DISABLED";
    FD1S3AX start_cnt_2121__i13 (.D(n10485), .CK(clkout_c), .Q(start_cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(391[18:27])
    defparam start_cnt_2121__i13.GSR = "DISABLED";
    AVG_SPEED_U9 AVG_SPEED_M3 (.\speed_avg_m3[0] (speed_avg_m3[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m3[0] (speed_m3[0]), .\speed_avg_m3[1] (speed_avg_m3[1]), 
            .\speed_m3[1] (speed_m3[1]), .\speed_avg_m3[2] (speed_avg_m3[2]), 
            .\speed_m3[2] (speed_m3[2]), .\speed_avg_m3[3] (speed_avg_m3[3]), 
            .\speed_m3[3] (speed_m3[3]), .\speed_avg_m3[4] (speed_avg_m3[4]), 
            .\speed_m3[4] (speed_m3[4]), .\speed_avg_m3[5] (speed_avg_m3[5]), 
            .\speed_m3[5] (speed_m3[5]), .\speed_avg_m3[6] (speed_avg_m3[6]), 
            .\speed_m3[6] (speed_m3[6]), .\speed_avg_m3[7] (speed_avg_m3[7]), 
            .\speed_m3[7] (speed_m3[7]), .\speed_avg_m3[8] (speed_avg_m3[8]), 
            .\speed_m3[8] (speed_m3[8]), .\speed_avg_m3[9] (speed_avg_m3[9]), 
            .\speed_m3[9] (speed_m3[9]), .\speed_avg_m3[10] (speed_avg_m3[10]), 
            .\speed_m3[10] (speed_m3[10]), .\speed_avg_m3[11] (speed_avg_m3[11]), 
            .\speed_m3[11] (speed_m3[11]), .\speed_avg_m3[12] (speed_avg_m3[12]), 
            .\speed_m3[12] (speed_m3[12]), .\speed_avg_m3[13] (speed_avg_m3[13]), 
            .\speed_m3[13] (speed_m3[13]), .\speed_avg_m3[14] (speed_avg_m3[14]), 
            .\speed_m3[14] (speed_m3[14]), .\speed_avg_m3[15] (speed_avg_m3[15]), 
            .\speed_m3[15] (speed_m3[15]), .\speed_avg_m3[16] (speed_avg_m3[16]), 
            .\speed_m3[16] (speed_m3[16]), .\speed_avg_m3[17] (speed_avg_m3[17]), 
            .\speed_m3[17] (speed_m3[17]), .\speed_avg_m3[18] (speed_avg_m3[18]), 
            .\speed_m3[18] (speed_m3[18]), .\speed_avg_m3[19] (speed_avg_m3[19]), 
            .\speed_m3[19] (speed_m3[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(367[17:26])
    AVG_SPEED_U10 AVG_SPEED_M2 (.\speed_avg_m2[0] (speed_avg_m2[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m2[0] (speed_m2[0]), .\speed_avg_m2[1] (speed_avg_m2[1]), 
            .\speed_m2[1] (speed_m2[1]), .\speed_avg_m2[2] (speed_avg_m2[2]), 
            .\speed_m2[2] (speed_m2[2]), .\speed_avg_m2[3] (speed_avg_m2[3]), 
            .\speed_m2[3] (speed_m2[3]), .\speed_avg_m2[4] (speed_avg_m2[4]), 
            .\speed_m2[4] (speed_m2[4]), .\speed_avg_m2[5] (speed_avg_m2[5]), 
            .\speed_m2[5] (speed_m2[5]), .\speed_avg_m2[6] (speed_avg_m2[6]), 
            .\speed_m2[6] (speed_m2[6]), .\speed_avg_m2[7] (speed_avg_m2[7]), 
            .\speed_m2[7] (speed_m2[7]), .\speed_avg_m2[8] (speed_avg_m2[8]), 
            .\speed_m2[8] (speed_m2[8]), .\speed_avg_m2[9] (speed_avg_m2[9]), 
            .\speed_m2[9] (speed_m2[9]), .\speed_avg_m2[10] (speed_avg_m2[10]), 
            .\speed_m2[10] (speed_m2[10]), .\speed_avg_m2[11] (speed_avg_m2[11]), 
            .\speed_m2[11] (speed_m2[11]), .\speed_avg_m2[12] (speed_avg_m2[12]), 
            .\speed_m2[12] (speed_m2[12]), .\speed_avg_m2[13] (speed_avg_m2[13]), 
            .\speed_m2[13] (speed_m2[13]), .\speed_avg_m2[14] (speed_avg_m2[14]), 
            .\speed_m2[14] (speed_m2[14]), .\speed_avg_m2[15] (speed_avg_m2[15]), 
            .\speed_m2[15] (speed_m2[15]), .\speed_avg_m2[16] (speed_avg_m2[16]), 
            .\speed_m2[16] (speed_m2[16]), .\speed_avg_m2[17] (speed_avg_m2[17]), 
            .\speed_m2[17] (speed_m2[17]), .\speed_avg_m2[18] (speed_avg_m2[18]), 
            .\speed_m2[18] (speed_m2[18]), .\speed_avg_m2[19] (speed_avg_m2[19]), 
            .\speed_m2[19] (speed_m2[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(364[17:26])
    AVG_SPEED_U11 AVG_SPEED_M1 (.\speed_avg_m1[0] (speed_avg_m1[0]), .clk_1mhz(clk_1mhz), 
            .\speed_m1[0] (speed_m1[0]), .\speed_avg_m1[1] (speed_avg_m1[1]), 
            .\speed_m1[1] (speed_m1[1]), .\speed_avg_m1[2] (speed_avg_m1[2]), 
            .\speed_m1[2] (speed_m1[2]), .\speed_avg_m1[3] (speed_avg_m1[3]), 
            .\speed_m1[3] (speed_m1[3]), .\speed_avg_m1[4] (speed_avg_m1[4]), 
            .\speed_m1[4] (speed_m1[4]), .\speed_avg_m1[5] (speed_avg_m1[5]), 
            .\speed_m1[5] (speed_m1[5]), .\speed_avg_m1[6] (speed_avg_m1[6]), 
            .\speed_m1[6] (speed_m1[6]), .\speed_avg_m1[7] (speed_avg_m1[7]), 
            .\speed_m1[7] (speed_m1[7]), .\speed_avg_m1[8] (speed_avg_m1[8]), 
            .\speed_m1[8] (speed_m1[8]), .\speed_avg_m1[9] (speed_avg_m1[9]), 
            .\speed_m1[9] (speed_m1[9]), .\speed_avg_m1[10] (speed_avg_m1[10]), 
            .\speed_m1[10] (speed_m1[10]), .\speed_avg_m1[11] (speed_avg_m1[11]), 
            .\speed_m1[11] (speed_m1[11]), .\speed_avg_m1[12] (speed_avg_m1[12]), 
            .\speed_m1[12] (speed_m1[12]), .\speed_avg_m1[13] (speed_avg_m1[13]), 
            .\speed_m1[13] (speed_m1[13]), .\speed_avg_m1[14] (speed_avg_m1[14]), 
            .\speed_m1[14] (speed_m1[14]), .\speed_avg_m1[15] (speed_avg_m1[15]), 
            .\speed_m1[15] (speed_m1[15]), .\speed_avg_m1[16] (speed_avg_m1[16]), 
            .\speed_m1[16] (speed_m1[16]), .\speed_avg_m1[17] (speed_avg_m1[17]), 
            .\speed_m1[17] (speed_m1[17]), .\speed_avg_m1[18] (speed_avg_m1[18]), 
            .\speed_m1[18] (speed_m1[18]), .\speed_avg_m1[19] (speed_avg_m1[19]), 
            .\speed_m1[19] (speed_m1[19]), .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(361[17:26])
    PWMGENERATOR_U1 PWM_I_M2 (.PWM_m2(PWM_m2), .pwm_clk(pwm_clk), .LED2_c(LED2_c), 
            .clkout_c_enable_362(clkout_c_enable_362), .PWMdut_m2({PWMdut_m2}), 
            .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(338[13:25])
    PWMGENERATOR_U0 PWM_I_M3 (.PWMdut_m3({PWMdut_m3}), .GND_net(GND_net), 
            .PWM_m3(PWM_m3), .pwm_clk(pwm_clk), .LED3_c(LED3_c), .clkout_c_enable_362(clkout_c_enable_362));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(348[13:25])
    PWMGENERATOR_U2 PWM_I_M1 (.PWMdut_m1({PWMdut_m1}), .GND_net(GND_net), 
            .PWM_m1(PWM_m1), .pwm_clk(pwm_clk), .LED1_c(LED1_c), .clkout_c_enable_362(clkout_c_enable_362));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(328[13:25])
    \PID(16000000,160000000,10000000)  PID_I (.speed_set_m2({speed_set_m2}), 
            .GND_net(GND_net), .clk_N_875(clk_N_875), .speed_set_m3({speed_set_m3}), 
            .\subOut_24__N_1369[0] (subOut_24__N_1369[0]), .speed_set_m1({speed_set_m1}), 
            .speed_set_m4({speed_set_m4}), .dir_m2(dir_m2), .dir_m3(dir_m3), 
            .dir_m1(dir_m1), .dir_m4(dir_m4), .\speed_avg_m3[12] (speed_avg_m3[12]), 
            .\speed_avg_m2[12] (speed_avg_m2[12]), .\speed_avg_m1[12] (speed_avg_m1[12]), 
            .\speed_avg_m1[9] (speed_avg_m1[9]), .\speed_avg_m1[8] (speed_avg_m1[8]), 
            .\speed_avg_m1[7] (speed_avg_m1[7]), .\speed_avg_m1[3] (speed_avg_m1[3]), 
            .\speed_avg_m1[19] (speed_avg_m1[19]), .\speed_avg_m2[19] (speed_avg_m2[19]), 
            .VCC_net(VCC_net), .\speed_avg_m1[18] (speed_avg_m1[18]), .\speed_avg_m2[18] (speed_avg_m2[18]), 
            .\speed_avg_m1[17] (speed_avg_m1[17]), .\speed_avg_m2[17] (speed_avg_m2[17]), 
            .\speed_avg_m1[16] (speed_avg_m1[16]), .\speed_avg_m2[16] (speed_avg_m2[16]), 
            .\speed_avg_m1[15] (speed_avg_m1[15]), .\speed_avg_m2[15] (speed_avg_m2[15]), 
            .\speed_avg_m1[14] (speed_avg_m1[14]), .\speed_avg_m2[14] (speed_avg_m2[14]), 
            .\speed_avg_m1[13] (speed_avg_m1[13]), .\speed_avg_m2[13] (speed_avg_m2[13]), 
            .\speed_avg_m1[11] (speed_avg_m1[11]), .\speed_avg_m2[11] (speed_avg_m2[11]), 
            .\speed_avg_m1[10] (speed_avg_m1[10]), .\speed_avg_m2[10] (speed_avg_m2[10]), 
            .\speed_avg_m1[6] (speed_avg_m1[6]), .\speed_avg_m2[6] (speed_avg_m2[6]), 
            .\speed_avg_m1[5] (speed_avg_m1[5]), .\speed_avg_m2[5] (speed_avg_m2[5]), 
            .\speed_avg_m1[4] (speed_avg_m1[4]), .\speed_avg_m2[4] (speed_avg_m2[4]), 
            .\speed_avg_m1[2] (speed_avg_m1[2]), .\speed_avg_m2[2] (speed_avg_m2[2]), 
            .\speed_avg_m3[9] (speed_avg_m3[9]), .\speed_avg_m2[9] (speed_avg_m2[9]), 
            .\speed_avg_m1[1] (speed_avg_m1[1]), .\speed_avg_m2[1] (speed_avg_m2[1]), 
            .\speed_avg_m1[0] (speed_avg_m1[0]), .\speed_avg_m2[0] (speed_avg_m2[0]), 
            .n19649(n19649), .\speed_avg_m3[8] (speed_avg_m3[8]), .\speed_avg_m2[8] (speed_avg_m2[8]), 
            .\speed_avg_m3[7] (speed_avg_m3[7]), .\speed_avg_m2[7] (speed_avg_m2[7]), 
            .\speed_avg_m3[3] (speed_avg_m3[3]), .\speed_avg_m2[3] (speed_avg_m2[3]), 
            .\speed_avg_m4[19] (speed_avg_m4[19]), .\speed_avg_m3[19] (speed_avg_m3[19]), 
            .\speed_avg_m4[18] (speed_avg_m4[18]), .\speed_avg_m3[18] (speed_avg_m3[18]), 
            .\speed_avg_m4[17] (speed_avg_m4[17]), .\speed_avg_m3[17] (speed_avg_m3[17]), 
            .\speed_avg_m4[16] (speed_avg_m4[16]), .\speed_avg_m3[16] (speed_avg_m3[16]), 
            .\speed_avg_m4[15] (speed_avg_m4[15]), .\speed_avg_m3[15] (speed_avg_m3[15]), 
            .\speed_avg_m4[14] (speed_avg_m4[14]), .\speed_avg_m3[14] (speed_avg_m3[14]), 
            .\speed_avg_m4[13] (speed_avg_m4[13]), .\speed_avg_m3[13] (speed_avg_m3[13]), 
            .\speed_avg_m4[11] (speed_avg_m4[11]), .\speed_avg_m3[11] (speed_avg_m3[11]), 
            .\speed_avg_m4[10] (speed_avg_m4[10]), .\speed_avg_m3[10] (speed_avg_m3[10]), 
            .\subOut_24__N_1369[1] (subOut_24__N_1369[1]), .\subOut_24__N_1369[2] (subOut_24__N_1369[2]), 
            .\subOut_24__N_1369[3] (subOut_24__N_1369[3]), .\subOut_24__N_1369[4] (subOut_24__N_1369[4]), 
            .\subOut_24__N_1369[5] (subOut_24__N_1369[5]), .\subOut_24__N_1369[6] (subOut_24__N_1369[6]), 
            .\subOut_24__N_1369[7] (subOut_24__N_1369[7]), .\subOut_24__N_1369[8] (subOut_24__N_1369[8]), 
            .\subOut_24__N_1369[9] (subOut_24__N_1369[9]), .\subOut_24__N_1369[10] (subOut_24__N_1369[10]), 
            .\subOut_24__N_1369[11] (subOut_24__N_1369[11]), .\subOut_24__N_1369[12] (subOut_24__N_1369[12]), 
            .\subOut_24__N_1369[13] (subOut_24__N_1369[13]), .\subOut_24__N_1369[14] (subOut_24__N_1369[14]), 
            .\subOut_24__N_1369[15] (subOut_24__N_1369[15]), .\subOut_24__N_1369[16] (subOut_24__N_1369[16]), 
            .\subOut_24__N_1369[17] (subOut_24__N_1369[17]), .\subOut_24__N_1369[18] (subOut_24__N_1369[18]), 
            .\subOut_24__N_1369[19] (subOut_24__N_1369[19]), .\subOut_24__N_1369[20] (subOut_24__N_1369[20]), 
            .\subOut_24__N_1369[21] (subOut_24__N_1369[21]), .\subOut_24__N_1369[24] (subOut_24__N_1369[24]), 
            .\speed_avg_m4[6] (speed_avg_m4[6]), .\speed_avg_m3[6] (speed_avg_m3[6]), 
            .\speed_avg_m4[5] (speed_avg_m4[5]), .\speed_avg_m3[5] (speed_avg_m3[5]), 
            .\speed_avg_m4[4] (speed_avg_m4[4]), .\speed_avg_m3[4] (speed_avg_m3[4]), 
            .\speed_avg_m4[2] (speed_avg_m4[2]), .\speed_avg_m3[2] (speed_avg_m3[2]), 
            .\speed_avg_m4[1] (speed_avg_m4[1]), .\speed_avg_m3[1] (speed_avg_m3[1]), 
            .\speed_avg_m4[0] (speed_avg_m4[0]), .\speed_avg_m3[0] (speed_avg_m3[0]), 
            .\speed_avg_m4[12] (speed_avg_m4[12]), .\speed_avg_m4[9] (speed_avg_m4[9]), 
            .\speed_avg_m4[8] (speed_avg_m4[8]), .\speed_avg_m4[7] (speed_avg_m4[7]), 
            .\speed_avg_m4[3] (speed_avg_m4[3]), .n22211(n22211), .PWMdut_m4({PWMdut_m4}), 
            .PWMdut_m3({PWMdut_m3}), .PWMdut_m2({PWMdut_m2}), .PWMdut_m1({PWMdut_m1}), 
            .n4510(n4510), .n4512(n4512), .n4511(n4511), .n4514(n4514), 
            .n4513(n4513), .n4516(n4516), .n4515(n4515), .n4518(n4518), 
            .n4517(n4517), .n4520(n4520), .n4519(n4519), .n4522(n4522), 
            .n4521(n4521), .n4524(n4524), .n4523(n4523), .n4526(n4526), 
            .n4525(n4525), .n4528(n4528), .n4527(n4527), .n4530(n4530), 
            .n4529(n4529), .n4531(n4531), .n4485(n4485), .n4484(n4484), 
            .n4487(n4487), .n4486(n4486), .n4489(n4489), .n4488(n4488), 
            .n4491(n4491), .n4490(n4490), .n4493(n4493), .n4492(n4492), 
            .n4495(n4495), .n4494(n4494), .n4497(n4497), .n4496(n4496), 
            .n4499(n4499), .n4498(n4498), .n4501(n4501), .n4500(n4500), 
            .n4503(n4503), .n4502(n4502), .n4505(n4505), .n4504(n4504), 
            .n4506(n4506));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(317[10:13])
    PWMGENERATOR PWM_I_M4 (.pwm_clk(pwm_clk), .PWM_m4(PWM_m4), .LED4_c(LED4_c), 
            .clkout_c_enable_362(clkout_c_enable_362), .PWMdut_m4({PWMdut_m4}), 
            .GND_net(GND_net));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(358[13:25])
    HALL HALL_I_M4 (.clk_1mhz(clk_1mhz), .\speed_m4[0] (speed_m4[0]), .hallsense_m4({hallsense_m4}), 
         .clkout_c_enable_266(clkout_c_enable_266), .clkout_c_enable_362(clkout_c_enable_362), 
         .H_A_m4_c(H_A_m4_c), .H_B_m4_c(H_B_m4_c), .H_C_m4_c(H_C_m4_c), 
         .\speed_m4[1] (speed_m4[1]), .\speed_m4[2] (speed_m4[2]), .\speed_m4[3] (speed_m4[3]), 
         .\speed_m4[4] (speed_m4[4]), .\speed_m4[5] (speed_m4[5]), .\speed_m4[6] (speed_m4[6]), 
         .\speed_m4[7] (speed_m4[7]), .\speed_m4[8] (speed_m4[8]), .\speed_m4[9] (speed_m4[9]), 
         .\speed_m4[10] (speed_m4[10]), .\speed_m4[11] (speed_m4[11]), .\speed_m4[12] (speed_m4[12]), 
         .\speed_m4[13] (speed_m4[13]), .\speed_m4[14] (speed_m4[14]), .\speed_m4[15] (speed_m4[15]), 
         .\speed_m4[16] (speed_m4[16]), .\speed_m4[17] (speed_m4[17]), .\speed_m4[18] (speed_m4[18]), 
         .\speed_m4[19] (speed_m4[19]), .GND_net(GND_net), .n22206(n22206));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(352[14:18])
    
endmodule
//
// Verilog Description of module CLKDIV
//

module CLKDIV (clk_N_875, clkout_c, clk_1mhz, pwm_clk, GND_net);
    output clk_N_875;
    input clkout_c;
    output clk_1mhz;
    output pwm_clk;
    input GND_net;
    
    wire clk_N_875 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    wire pi_clk /* synthesis is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(89[9:15])
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire mhz_buf, mhz_buf_N_68, pi_buf, pi_buf_N_69, pwm_buf, pwm_buf_N_67;
    wire [4:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(41[8:13])
    
    wire n14212;
    wire [4:0]n25;
    
    wire n19707, n14211, n15;
    wire [11:0]cntpi;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(42[8:13])
    
    wire n14, n21477;
    wire [8:0]n41;
    
    wire n18362, n18361, n18360, n18359;
    
    INV i17535 (.A(pi_clk), .Z(clk_N_875));
    FD1S3AX mhz_buf_29 (.D(mhz_buf_N_68), .CK(clkout_c), .Q(mhz_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=308, LSE_RLINE=308 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam mhz_buf_29.GSR = "DISABLED";
    FD1S3AX pi_buf_30 (.D(pi_buf_N_69), .CK(clkout_c), .Q(pi_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=308, LSE_RLINE=308 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pi_buf_30.GSR = "DISABLED";
    FD1S3AX pwm_buf_32 (.D(pwm_buf_N_67), .CK(clkout_c), .Q(pwm_buf)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=308, LSE_RLINE=308 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pwm_buf_32.GSR = "DISABLED";
    FD1S3AX clk_1mhz_33 (.D(mhz_buf), .CK(clkout_c), .Q(clk_1mhz)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=308, LSE_RLINE=308 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam clk_1mhz_33.GSR = "DISABLED";
    FD1S3AX pwm_clk_34 (.D(pwm_buf), .CK(clkout_c), .Q(pwm_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=308, LSE_RLINE=308 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pwm_clk_34.GSR = "DISABLED";
    FD1S3AX pi_clk_35 (.D(pi_buf), .CK(clkout_c), .Q(pi_clk)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=20, LSE_LLINE=308, LSE_RLINE=308 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(55[1] 79[8])
    defparam pi_clk_35.GSR = "DISABLED";
    FD1S3IX count_2122__i0 (.D(n25[0]), .CK(clkout_c), .CD(n14212), .Q(count[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2122__i0.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(mhz_buf), .B(n14212), .Z(mhz_buf_N_68)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    LUT4 i17186_4_lut (.A(count[2]), .B(count[0]), .C(count[3]), .D(n19707), 
         .Z(n14212)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(61[5:15])
    defparam i17186_4_lut.init = 16'h0400;
    LUT4 i16256_2_lut (.A(count[4]), .B(count[1]), .Z(n19707)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16256_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_190 (.A(pi_buf), .B(n14211), .Z(pi_buf_N_69)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_190.init = 16'h6666;
    LUT4 i17183_4_lut (.A(n15), .B(cntpi[6]), .C(n14), .D(cntpi[4]), 
         .Z(n14211)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(66[5:16])
    defparam i17183_4_lut.init = 16'h0400;
    LUT4 i6_4_lut (.A(cntpi[7]), .B(cntpi[0]), .C(cntpi[1]), .D(cntpi[5]), 
         .Z(n15)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'hbfff;
    LUT4 i15175_3_lut_4_lut (.A(count[2]), .B(n21477), .C(count[3]), .D(count[4]), 
         .Z(n25[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15175_3_lut_4_lut.init = 16'h7f80;
    LUT4 i5_3_lut (.A(cntpi[3]), .B(cntpi[8]), .C(cntpi[2]), .Z(n14)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i5_3_lut.init = 16'hf7f7;
    LUT4 pwm_buf_I_0_1_lut (.A(pwm_buf), .Z(pwm_buf_N_67)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(73[14:25])
    defparam pwm_buf_I_0_1_lut.init = 16'h5555;
    LUT4 i15152_1_lut (.A(count[0]), .Z(n25[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15152_1_lut.init = 16'h5555;
    LUT4 i15157_2_lut_rep_376 (.A(count[1]), .B(count[0]), .Z(n21477)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15157_2_lut_rep_376.init = 16'h8888;
    LUT4 i15161_2_lut_3_lut (.A(count[1]), .B(count[0]), .C(count[2]), 
         .Z(n25[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15161_2_lut_3_lut.init = 16'h7878;
    LUT4 i15168_2_lut_3_lut_4_lut (.A(count[1]), .B(count[0]), .C(count[3]), 
         .D(count[2]), .Z(n25[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15168_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i15154_2_lut (.A(count[1]), .B(count[0]), .Z(n25[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam i15154_2_lut.init = 16'h6666;
    FD1S3IX cntpi_2123_2124__i2 (.D(n41[1]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i2.GSR = "DISABLED";
    FD1S3IX cntpi_2123_2124__i1 (.D(n41[0]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i1.GSR = "DISABLED";
    CCU2D cntpi_2123_2124_add_4_9 (.A0(cntpi[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18362), .S0(n41[7]), .S1(n41[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124_add_4_9.INIT0 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_9.INIT1 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_9.INJECT1_0 = "NO";
    defparam cntpi_2123_2124_add_4_9.INJECT1_1 = "NO";
    CCU2D cntpi_2123_2124_add_4_7 (.A0(cntpi[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18361), .COUT(n18362), .S0(n41[5]), .S1(n41[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124_add_4_7.INIT0 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_7.INIT1 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_7.INJECT1_0 = "NO";
    defparam cntpi_2123_2124_add_4_7.INJECT1_1 = "NO";
    CCU2D cntpi_2123_2124_add_4_5 (.A0(cntpi[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18360), .COUT(n18361), .S0(n41[3]), .S1(n41[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124_add_4_5.INIT0 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_5.INIT1 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_5.INJECT1_0 = "NO";
    defparam cntpi_2123_2124_add_4_5.INJECT1_1 = "NO";
    CCU2D cntpi_2123_2124_add_4_3 (.A0(cntpi[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18359), .COUT(n18360), .S0(n41[1]), .S1(n41[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124_add_4_3.INIT0 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_3.INIT1 = 16'hfaaa;
    defparam cntpi_2123_2124_add_4_3.INJECT1_0 = "NO";
    defparam cntpi_2123_2124_add_4_3.INJECT1_1 = "NO";
    CCU2D cntpi_2123_2124_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cntpi[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18359), .S1(n41[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124_add_4_1.INIT0 = 16'hF000;
    defparam cntpi_2123_2124_add_4_1.INIT1 = 16'h0555;
    defparam cntpi_2123_2124_add_4_1.INJECT1_0 = "NO";
    defparam cntpi_2123_2124_add_4_1.INJECT1_1 = "NO";
    FD1S3IX cntpi_2123_2124__i3 (.D(n41[2]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i3.GSR = "DISABLED";
    FD1S3IX cntpi_2123_2124__i4 (.D(n41[3]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i4.GSR = "DISABLED";
    FD1S3IX cntpi_2123_2124__i5 (.D(n41[4]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i5.GSR = "DISABLED";
    FD1S3IX cntpi_2123_2124__i6 (.D(n41[5]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i6.GSR = "DISABLED";
    FD1S3IX cntpi_2123_2124__i7 (.D(n41[6]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i7.GSR = "DISABLED";
    FD1S3IX cntpi_2123_2124__i8 (.D(n41[7]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i8.GSR = "DISABLED";
    FD1S3IX cntpi_2123_2124__i9 (.D(n41[8]), .CK(clkout_c), .CD(n14211), 
            .Q(cntpi[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(57[11:16])
    defparam cntpi_2123_2124__i9.GSR = "DISABLED";
    FD1S3IX count_2122__i1 (.D(n25[1]), .CK(clkout_c), .CD(n14212), .Q(count[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2122__i1.GSR = "DISABLED";
    FD1S3IX count_2122__i2 (.D(n25[2]), .CK(clkout_c), .CD(n14212), .Q(count[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2122__i2.GSR = "DISABLED";
    FD1S3IX count_2122__i3 (.D(n25[3]), .CK(clkout_c), .CD(n14212), .Q(count[3]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2122__i3.GSR = "DISABLED";
    FD1S3IX count_2122__i4 (.D(n25[4]), .CK(clkout_c), .CD(n14212), .Q(count[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/clockdivider.vhd(56[11:16])
    defparam count_2122__i4.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module HALL_U4
//

module HALL_U4 (clk_1mhz, \speed_m2[0] , hallsense_m2, rst, H_B_m2_c, 
            clkout_c_enable_266, H_A_m2_c, clkout_c_enable_362, H_C_m2_c, 
            \speed_m2[1] , \speed_m2[2] , \speed_m2[3] , \speed_m2[4] , 
            \speed_m2[5] , \speed_m2[6] , \speed_m2[7] , \speed_m2[8] , 
            \speed_m2[9] , \speed_m2[10] , \speed_m2[11] , \speed_m2[12] , 
            \speed_m2[13] , \speed_m2[14] , \speed_m2[15] , \speed_m2[16] , 
            \speed_m2[17] , \speed_m2[18] , \speed_m2[19] , GND_net, 
            n22206);
    input clk_1mhz;
    output \speed_m2[0] ;
    output [2:0]hallsense_m2;
    input rst;
    input H_B_m2_c;
    input clkout_c_enable_266;
    input H_A_m2_c;
    input clkout_c_enable_362;
    input H_C_m2_c;
    output \speed_m2[1] ;
    output \speed_m2[2] ;
    output \speed_m2[3] ;
    output \speed_m2[4] ;
    output \speed_m2[5] ;
    output \speed_m2[6] ;
    output \speed_m2[7] ;
    output \speed_m2[8] ;
    output \speed_m2[9] ;
    output \speed_m2[10] ;
    output \speed_m2[11] ;
    output \speed_m2[12] ;
    output \speed_m2[13] ;
    output \speed_m2[14] ;
    output \speed_m2[15] ;
    output \speed_m2[16] ;
    output \speed_m2[17] ;
    output \speed_m2[18] ;
    output \speed_m2[19] ;
    input GND_net;
    input n22206;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_50;
    wire [19:0]count_19__N_2069;
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21460, n21416, n4, stable_counting;
    wire [19:0]speedt_19__N_2049;
    
    wire hall3_lat;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4621, hall2_lat, hall1_lat, hall3_old, hall1_old, hall2_old, 
        n11577, n11575, stable_counting_N_2131, n13, n12, n19873, 
        n19877, n19875, n19731, n19657, n21426, n19574, n21412;
    wire [6:0]n63;
    
    wire n4_adj_2426, n18858, n19789, clk_1mhz_enable_186, n25, n26, 
        n22, n19859, n19857, n24, n18, n21425, n21486, n21461, 
        n21441, n14446, n18293, n18292, n18291, n18290, n18289, 
        n18288, n18287, n18286, n18285, n18284;
    
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2069[0]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    LUT4 i2485_2_lut_rep_315_3_lut_4_lut (.A(stable_count[3]), .B(n21460), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21416)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2485_2_lut_rep_315_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21460), .C(stable_count[0]), 
         .D(stable_count[4]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h7f8f;
    FD1P3AX speed__i1 (.D(speedt_19__N_2049[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_19__N_2069[0]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m2_c), .SP(rst), .CK(clk_1mhz), .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(H_A_m2_c), .SP(clkout_c_enable_266), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m2_c), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2069[1]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2069[17]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2069[16]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2069[15]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2069[14]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2069[13]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2069[12]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2069[11]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2069[10]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2069[9]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2069[8]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2069[7]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2069[6]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2069[5]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2069[4]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2069[19]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2069[3]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2069[18]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2069[2]), .SP(clk_1mhz_enable_50), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2049[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2049[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2049[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2049[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2049[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2049[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2049[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2049[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2049[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2049[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2049[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2049[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2049[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i11564_4_lut (.A(n11577), .B(n11575), .C(stable_counting), .D(stable_counting_N_2131), 
         .Z(clk_1mhz_enable_50)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11564_4_lut.init = 16'hcaea;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2049[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2049[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7_4_lut (.A(n13), .B(count[2]), .C(n12), .D(count[10]), .Z(n11577)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[9]), .B(count[3]), .C(count[8]), .D(count[13]), 
         .Z(n13)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2049[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2049[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4_4_lut (.A(count[0]), .B(n19873), .C(n19877), .D(n19875), 
         .Z(n12)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h0002;
    LUT4 i16421_4_lut (.A(count[7]), .B(count[14]), .C(count[6]), .D(n19731), 
         .Z(n19873)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16421_4_lut.init = 16'hfffe;
    LUT4 i16425_4_lut (.A(count[18]), .B(count[19]), .C(count[11]), .D(count[16]), 
         .Z(n19877)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16425_4_lut.init = 16'hfffe;
    LUT4 i16423_4_lut (.A(count[4]), .B(count[5]), .C(count[17]), .D(count[1]), 
         .Z(n19875)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16423_4_lut.init = 16'hfffe;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2049[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16280_2_lut (.A(count[12]), .B(count[15]), .Z(n19731)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16280_2_lut.init = 16'heeee;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2049[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11577), .B(n11575), .C(count_19__N_2069[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2049[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_4_lut (.A(n19657), .B(stable_count[0]), .C(n21426), .D(n19574), 
         .Z(n11575)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    LUT4 i2_4_lut_adj_187 (.A(n19657), .B(n21412), .C(n63[2]), .D(n4), 
         .Z(stable_counting_N_2131)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i2_4_lut_adj_187.init = 16'h0002;
    LUT4 i1_4_lut (.A(hall2_old), .B(hall1_old), .C(hall2_lat), .D(hall1_lat), 
         .Z(n4_adj_2426)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i2457_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2457_2_lut.init = 16'h6666;
    FD1P3AX speed__i2 (.D(speedt_19__N_2049[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2049[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2049[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2049[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2049[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2049[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2049[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2049[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m2[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2049[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2049[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2049[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2049[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2049[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2049[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2049[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2049[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2049[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2049[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2049[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m2[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i2292_2_lut (.A(stable_counting), .B(stable_counting_N_2131), .Z(n4621)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2292_2_lut.init = 16'h8888;
    FD1S3IX count__i1 (.D(count_19__N_2069[1]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2069[2]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2069[3]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2069[4]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2069[5]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2069[6]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2069[7]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2069[8]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2069[9]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2069[10]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2069[11]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2069[12]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2069[13]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2069[14]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2069[15]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2069[16]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2069[17]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2069[18]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2069[19]), .CK(clk_1mhz), .CD(n4621), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n21416), .B(n63[6]), .C(n63[3]), .D(n63[2]), 
         .Z(n19574)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i17259_4_lut (.A(n18858), .B(n19789), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_186)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17259_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_188 (.A(n25), .B(count[0]), .C(n26), .D(count[10]), 
         .Z(n18858)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i1_4_lut_adj_188.init = 16'hfbff;
    LUT4 i16338_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19789)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16338_4_lut.init = 16'h7bde;
    LUT4 i11_4_lut (.A(count[1]), .B(n22), .C(n19859), .D(n19857), .Z(n25)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i11_4_lut.init = 16'hefff;
    LUT4 i12_4_lut (.A(count[5]), .B(n24), .C(n18), .D(count[19]), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[17]), .B(count[16]), .C(count[18]), .D(count[15]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i16407_2_lut (.A(count[8]), .B(count[13]), .Z(n19859)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16407_2_lut.init = 16'h8888;
    LUT4 i16405_3_lut (.A(count[2]), .B(count[3]), .C(count[9]), .Z(n19857)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16405_3_lut.init = 16'h8080;
    LUT4 i10_4_lut (.A(count[11]), .B(count[6]), .C(count[7]), .D(count[14]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[4]), .B(count[12]), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_rep_311_4_lut (.A(stable_count[5]), .B(n21425), .C(n63[3]), 
         .D(n63[6]), .Z(n21412)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_311_4_lut.init = 16'hfff6;
    LUT4 i2455_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2455_1_lut.init = 16'h5555;
    LUT4 i2480_2_lut_rep_324_3_lut_4_lut (.A(stable_count[2]), .B(n21486), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21425)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2480_2_lut_rep_324_3_lut_4_lut.init = 16'h8000;
    LUT4 i2478_2_lut_rep_325_3_lut_4_lut (.A(stable_count[2]), .B(n21486), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21426)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2478_2_lut_rep_325_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2_3_lut_rep_360 (.A(hall3_old), .B(n4_adj_2426), .C(hall3_lat), 
         .Z(n21461)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_360.init = 16'hdede;
    LUT4 i1_2_lut_4_lut_adj_189 (.A(hall3_old), .B(n4_adj_2426), .C(hall3_lat), 
         .D(n63[1]), .Z(n19657)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_189.init = 16'h2100;
    LUT4 i2492_3_lut_4_lut (.A(stable_count[4]), .B(n21441), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2492_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2459_2_lut_rep_385 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21486)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2459_2_lut_rep_385.init = 16'h8888;
    LUT4 i2464_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2464_2_lut_3_lut.init = 16'h7878;
    LUT4 i16413_3_lut (.A(n21461), .B(stable_counting), .C(stable_counting_N_2131), 
         .Z(n14446)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16413_3_lut.init = 16'hc8c8;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21416), .SP(stable_counting), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21426), .SP(stable_counting), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    LUT4 i2466_2_lut_rep_359_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21460)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2466_2_lut_rep_359_3_lut.init = 16'h8080;
    LUT4 i2473_2_lut_rep_340_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21441)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2473_2_lut_rep_340_3_lut_4_lut.init = 16'h8000;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18293), 
          .S0(count_19__N_2069[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    LUT4 i2471_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2471_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18292), .COUT(n18293), .S0(count_19__N_2069[17]), .S1(count_19__N_2069[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18291), .COUT(n18292), .S0(count_19__N_2069[15]), .S1(count_19__N_2069[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18290), .COUT(n18291), .S0(count_19__N_2069[13]), .S1(count_19__N_2069[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18289), .COUT(n18290), .S0(count_19__N_2069[11]), .S1(count_19__N_2069[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18288), .COUT(n18289), .S0(count_19__N_2069[9]), .S1(count_19__N_2069[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18287), 
          .COUT(n18288), .S0(count_19__N_2069[7]), .S1(count_19__N_2069[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    FD1P3IX stable_counting_62 (.D(n22206), .SP(clk_1mhz_enable_186), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18286), 
          .COUT(n18287), .S0(count_19__N_2069[5]), .S1(count_19__N_2069[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18285), 
          .COUT(n18286), .S0(count_19__N_2069[3]), .S1(count_19__N_2069[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14446), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=332, LSE_RLINE=332 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18284), 
          .COUT(n18285), .S0(count_19__N_2069[1]), .S1(count_19__N_2069[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18284), 
          .S1(count_19__N_2069[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module COMMUTATION_U7
//

module COMMUTATION_U7 (MB_m2_c_0, clkout_c, MC_m2_c_0, n21487, dir_m2, 
            hallsense_m2, MA_m2_c_1, n21453, PWM_m2, MC_m2_c_1, n3037, 
            MB_m2_c_1, n3003, LED2_c, enable_m2, MA_m2_c_0, n14200);
    output MB_m2_c_0;
    input clkout_c;
    output MC_m2_c_0;
    output n21487;
    input dir_m2;
    input [2:0]hallsense_m2;
    output MA_m2_c_1;
    input n21453;
    input PWM_m2;
    output MC_m2_c_1;
    input n3037;
    output MB_m2_c_1;
    input n3003;
    input LED2_c;
    input enable_m2;
    output MA_m2_c_0;
    input n14200;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire [1:0]MospairB_1__N_2141;
    wire [1:0]MospairC_1__N_2143;
    
    wire n21502, n8, n21263, n16065;
    
    FD1S3AX MospairB_i1 (.D(MospairB_1__N_2141[0]), .CK(clkout_c), .Q(MB_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3AX MospairC_i1 (.D(MospairC_1__N_2143[0]), .CK(clkout_c), .Q(MC_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i1.GSR = "DISABLED";
    LUT4 n21487_bdd_4_lut (.A(n21487), .B(dir_m2), .C(hallsense_m2[2]), 
         .D(hallsense_m2[0]), .Z(n21502)) /* synthesis lut_function=(!((B ((D)+!C)+!B (C+!(D)))+!A)) */ ;
    defparam n21487_bdd_4_lut.init = 16'h0280;
    LUT4 i21_4_lut (.A(hallsense_m2[0]), .B(n21487), .C(hallsense_m2[1]), 
         .D(dir_m2), .Z(n8)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i21_4_lut.init = 16'h400a;
    FD1S3IX MospairA_i2 (.D(n21502), .CK(clkout_c), .CD(n21453), .Q(MA_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i2.GSR = "DISABLED";
    LUT4 PWM_m2_bdd_4_lut (.A(PWM_m2), .B(hallsense_m2[1]), .C(hallsense_m2[2]), 
         .D(dir_m2), .Z(n21263)) /* synthesis lut_function=((B (C+(D))+!B !(C (D)))+!A) */ ;
    defparam PWM_m2_bdd_4_lut.init = 16'hdff7;
    FD1S3IX MospairC_i2 (.D(n21487), .CK(clkout_c), .CD(n3037), .Q(MC_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n21487), .CK(clkout_c), .CD(n3003), .Q(MB_m2_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i17161_2_lut_rep_386 (.A(LED2_c), .B(enable_m2), .Z(n21487)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17161_2_lut_rep_386.init = 16'h4444;
    FD1S3JX MospairA_i1 (.D(n16065), .CK(clkout_c), .PD(n14200), .Q(MA_m2_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=335, LSE_RLINE=335 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i1.GSR = "DISABLED";
    LUT4 i17230_3_lut_4_lut (.A(LED2_c), .B(enable_m2), .C(n8), .D(PWM_m2), 
         .Z(MospairC_1__N_2143[0])) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17230_3_lut_4_lut.init = 16'h0444;
    LUT4 i17253_2_lut_3_lut (.A(LED2_c), .B(enable_m2), .C(PWM_m2), .Z(n16065)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17253_2_lut_3_lut.init = 16'h0404;
    LUT4 gnd_bdd_2_lut_17329_3_lut (.A(LED2_c), .B(enable_m2), .C(n21263), 
         .Z(MospairB_1__N_2141[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam gnd_bdd_2_lut_17329_3_lut.init = 16'h4040;
    
endmodule
//
// Verilog Description of module COMMUTATION_U8
//

module COMMUTATION_U8 (n21476, dir_m1, hallsense_m1, MA_m1_c_0, clkout_c, 
            n14195, MB_m1_c_0, MC_m1_c_0, MA_m1_c_1, n21451, LED1_c, 
            enable_m1, PWM_m1, MC_m1_c_1, n2935, MB_m1_c_1, n2901);
    output n21476;
    input dir_m1;
    input [2:0]hallsense_m1;
    output MA_m1_c_0;
    input clkout_c;
    input n14195;
    output MB_m1_c_0;
    output MC_m1_c_0;
    output MA_m1_c_1;
    input n21451;
    input LED1_c;
    input enable_m1;
    input PWM_m1;
    output MC_m1_c_1;
    input n2935;
    output MB_m1_c_1;
    input n2901;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire n21503, n16107;
    wire [1:0]MospairB_1__N_2141;
    wire [1:0]MospairC_1__N_2143;
    
    wire n8, n21321;
    
    LUT4 n21476_bdd_4_lut (.A(n21476), .B(dir_m1), .C(hallsense_m1[2]), 
         .D(hallsense_m1[0]), .Z(n21503)) /* synthesis lut_function=(!((B ((D)+!C)+!B (C+!(D)))+!A)) */ ;
    defparam n21476_bdd_4_lut.init = 16'h0280;
    FD1S3JX MospairA_i1 (.D(n16107), .CK(clkout_c), .PD(n14195), .Q(MA_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3AX MospairB_i1 (.D(MospairB_1__N_2141[0]), .CK(clkout_c), .Q(MB_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3AX MospairC_i1 (.D(MospairC_1__N_2143[0]), .CK(clkout_c), .Q(MC_m1_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i1.GSR = "DISABLED";
    LUT4 i21_4_lut (.A(hallsense_m1[0]), .B(n21476), .C(hallsense_m1[1]), 
         .D(dir_m1), .Z(n8)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i21_4_lut.init = 16'h400a;
    FD1S3IX MospairA_i2 (.D(n21503), .CK(clkout_c), .CD(n21451), .Q(MA_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i2.GSR = "DISABLED";
    LUT4 i17152_2_lut_rep_375 (.A(LED1_c), .B(enable_m1), .Z(n21476)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17152_2_lut_rep_375.init = 16'h4444;
    LUT4 i17255_2_lut_3_lut (.A(LED1_c), .B(enable_m1), .C(PWM_m1), .Z(n16107)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17255_2_lut_3_lut.init = 16'h0404;
    LUT4 i17134_3_lut_4_lut (.A(LED1_c), .B(enable_m1), .C(n8), .D(PWM_m1), 
         .Z(MospairC_1__N_2143[0])) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17134_3_lut_4_lut.init = 16'h0444;
    LUT4 gnd_bdd_2_lut_17332_3_lut (.A(LED1_c), .B(enable_m1), .C(n21321), 
         .Z(MospairB_1__N_2141[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam gnd_bdd_2_lut_17332_3_lut.init = 16'h4040;
    LUT4 PWM_m1_bdd_4_lut (.A(PWM_m1), .B(hallsense_m1[1]), .C(hallsense_m1[2]), 
         .D(dir_m1), .Z(n21321)) /* synthesis lut_function=((B (C+(D))+!B !(C (D)))+!A) */ ;
    defparam PWM_m1_bdd_4_lut.init = 16'hdff7;
    FD1S3IX MospairC_i2 (.D(n21476), .CK(clkout_c), .CD(n2935), .Q(MC_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n21476), .CK(clkout_c), .CD(n2901), .Q(MB_m1_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=325, LSE_RLINE=325 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module HALL_U5
//

module HALL_U5 (clk_1mhz, GND_net, \speed_m1[0] , hallsense_m1, clkout_c_enable_362, 
            clkout_c_enable_266, HALL_A_OUT_c_c, HALL_B_OUT_c_c, HALL_C_OUT_c_c, 
            \speed_m1[1] , \speed_m1[2] , \speed_m1[3] , \speed_m1[4] , 
            \speed_m1[5] , \speed_m1[6] , \speed_m1[7] , \speed_m1[8] , 
            \speed_m1[9] , \speed_m1[10] , \speed_m1[11] , \speed_m1[12] , 
            \speed_m1[13] , \speed_m1[14] , \speed_m1[15] , \speed_m1[16] , 
            \speed_m1[17] , \speed_m1[18] , \speed_m1[19] , n22206);
    input clk_1mhz;
    input GND_net;
    output \speed_m1[0] ;
    output [2:0]hallsense_m1;
    input clkout_c_enable_362;
    input clkout_c_enable_266;
    input HALL_A_OUT_c_c;
    input HALL_B_OUT_c_c;
    input HALL_C_OUT_c_c;
    output \speed_m1[1] ;
    output \speed_m1[2] ;
    output \speed_m1[3] ;
    output \speed_m1[4] ;
    output \speed_m1[5] ;
    output \speed_m1[6] ;
    output \speed_m1[7] ;
    output \speed_m1[8] ;
    output \speed_m1[9] ;
    output \speed_m1[10] ;
    output \speed_m1[11] ;
    output \speed_m1[12] ;
    output \speed_m1[13] ;
    output \speed_m1[14] ;
    output \speed_m1[15] ;
    output \speed_m1[16] ;
    output \speed_m1[17] ;
    output \speed_m1[18] ;
    output \speed_m1[19] ;
    input n22206;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire n21457, n4;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_69;
    wire [19:0]count_19__N_2069;
    
    wire n18283;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n18282, n18281, stable_counting;
    wire [19:0]speedt_19__N_2049;
    
    wire hall3_lat, n18280, n18279, n18278, n18277, n18276, n4616, 
        n18275;
    wire [6:0]n63;
    
    wire hall1_old, hall1_lat, hall2_old, hall2_lat, hall3_old, n18274, 
        n4_adj_2425, n21450, n19642, n11582, n11580, stable_counting_N_2131, 
        n19586, n19775, n19909, n19889, n19885, n19781, n21423, 
        n19571, n21411, n21414, n21419, n18854, n19801, clk_1mhz_enable_185, 
        n19, n24, n20, n22, n16, n21439, n21482, n12, n14472;
    
    LUT4 i1_2_lut_3_lut_4_lut (.A(stable_count[3]), .B(n21457), .C(stable_count[0]), 
         .D(stable_count[4]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h7f8f;
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2069[0]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18283), 
          .S0(count_19__N_2069[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18282), .COUT(n18283), .S0(count_19__N_2069[17]), .S1(count_19__N_2069[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18281), .COUT(n18282), .S0(count_19__N_2069[15]), .S1(count_19__N_2069[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    FD1P3AX speed__i1 (.D(speedt_19__N_2049[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18280), .COUT(n18281), .S0(count_19__N_2069[13]), .S1(count_19__N_2069[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18279), .COUT(n18280), .S0(count_19__N_2069[11]), .S1(count_19__N_2069[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18278), .COUT(n18279), .S0(count_19__N_2069[9]), .S1(count_19__N_2069[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18277), 
          .COUT(n18278), .S0(count_19__N_2069[7]), .S1(count_19__N_2069[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18276), 
          .COUT(n18277), .S0(count_19__N_2069[5]), .S1(count_19__N_2069[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    FD1S3IX count__i0 (.D(count_19__N_2069[0]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18275), 
          .COUT(n18276), .S0(count_19__N_2069[3]), .S1(count_19__N_2069[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    LUT4 i2405_1_lut (.A(stable_count[0]), .Z(n63[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2405_1_lut.init = 16'h5555;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_266), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    FD1P3AX hall1_lat_57 (.D(HALL_A_OUT_c_c), .SP(clkout_c_enable_266), 
            .CK(clk_1mhz), .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(HALL_B_OUT_c_c), .SP(clkout_c_enable_266), 
            .CK(clk_1mhz), .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(HALL_C_OUT_c_c), .SP(clkout_c_enable_266), 
            .CK(clk_1mhz), .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18274), 
          .COUT(n18275), .S0(count_19__N_2069[1]), .S1(count_19__N_2069[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18274), 
          .S1(count_19__N_2069[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_349 (.A(hall3_old), .B(n4_adj_2425), .C(hall3_lat), 
         .Z(n21450)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_349.init = 16'hdede;
    LUT4 i1_2_lut_4_lut (.A(hall3_old), .B(n4_adj_2425), .C(hall3_lat), 
         .D(n63[1]), .Z(n19642)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h2100;
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2069[19]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2069[18]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2069[17]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2069[16]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2069[15]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2069[14]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2069[13]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2069[12]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2069[11]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2069[10]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2069[9]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2069[8]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2069[7]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2069[6]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2069[5]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2069[4]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2069[3]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2069[2]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2069[1]), .SP(clk_1mhz_enable_69), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2049[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2049[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2049[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2049[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2049[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2049[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2049[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2049[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2049[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i11562_4_lut (.A(n11582), .B(n11580), .C(stable_counting), .D(stable_counting_N_2131), 
         .Z(clk_1mhz_enable_69)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11562_4_lut.init = 16'hcaea;
    LUT4 i1_4_lut (.A(n19586), .B(n19775), .C(n19909), .D(n19889), .Z(n11582)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0002;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2049[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2049[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16324_2_lut (.A(count[18]), .B(count[1]), .Z(n19775)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16324_2_lut.init = 16'heeee;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2049[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2049[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2049[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX speed__i2 (.D(speedt_19__N_2049[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2049[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2049[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2049[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2049[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2049[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2049[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2049[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m1[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2049[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2049[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2049[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2049[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2049[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2049[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2049[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2049[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2049[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2049[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2049[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m1[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i16457_4_lut (.A(count[5]), .B(n19885), .C(n19781), .D(count[12]), 
         .Z(n19909)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16457_4_lut.init = 16'hfffe;
    LUT4 i16437_3_lut (.A(count[15]), .B(count[7]), .C(count[16]), .Z(n19889)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16437_3_lut.init = 16'hfefe;
    LUT4 i16433_4_lut (.A(count[11]), .B(count[17]), .C(count[4]), .D(count[6]), 
         .Z(n19885)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16433_4_lut.init = 16'hfffe;
    LUT4 i16330_2_lut (.A(count[19]), .B(count[14]), .Z(n19781)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16330_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(n21423), .B(stable_count[0]), .C(n19571), .D(n19642), 
         .Z(n11580)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i1_4_lut_adj_183 (.A(n63[2]), .B(n19642), .C(n21411), .D(n4), 
         .Z(stable_counting_N_2131)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_183.init = 16'h0004;
    LUT4 i2289_2_lut (.A(stable_counting), .B(stable_counting_N_2131), .Z(n4616)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2289_2_lut.init = 16'h8888;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2049[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2049[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2049[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX count__i1 (.D(count_19__N_2069[1]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2069[2]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2069[3]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2069[4]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2069[5]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2069[6]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2069[7]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2069[8]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2069[9]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2069[10]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2069[11]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2069[12]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2069[13]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2069[14]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2069[15]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2069[16]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2069[17]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2069[18]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2069[19]), .CK(clk_1mhz), .CD(n4616), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2049[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2049[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11582), .B(n11580), .C(count_19__N_2069[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2049[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_184 (.A(n21414), .B(n63[6]), .C(n63[3]), .D(n63[2]), 
         .Z(n19571)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_2_lut_4_lut_adj_184.init = 16'hfffe;
    LUT4 i2_3_lut_rep_310_4_lut (.A(stable_count[5]), .B(n21419), .C(n63[3]), 
         .D(n63[6]), .Z(n21411)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_310_4_lut.init = 16'hfff6;
    LUT4 i17261_4_lut (.A(n18854), .B(n19801), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_185)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17261_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_185 (.A(n19), .B(n19586), .C(n24), .D(n20), .Z(n18854)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i1_4_lut_adj_185.init = 16'hfffb;
    LUT4 i16349_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19801)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16349_4_lut.init = 16'h7bde;
    LUT4 i6_2_lut (.A(count[17]), .B(count[12]), .Z(n19)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i11_4_lut (.A(count[5]), .B(n22), .C(n16), .D(count[16]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut (.A(count[14]), .B(count[19]), .C(count[11]), .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i9_4_lut (.A(count[15]), .B(count[18]), .C(count[1]), .D(count[4]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(count[6]), .B(count[7]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i2442_3_lut_4_lut (.A(stable_count[4]), .B(n21439), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2442_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2430_2_lut_rep_318_3_lut_4_lut (.A(stable_count[2]), .B(n21482), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21419)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2430_2_lut_rep_318_3_lut_4_lut.init = 16'h8000;
    LUT4 i2428_2_lut_rep_322_3_lut_4_lut (.A(stable_count[2]), .B(n21482), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21423)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2428_2_lut_rep_322_3_lut_4_lut.init = 16'h78f0;
    LUT4 i6_4_lut (.A(count[0]), .B(n12), .C(count[9]), .D(count[8]), 
         .Z(n19586)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[3]), .B(count[2]), .C(count[13]), .D(count[10]), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i16415_3_lut (.A(n21450), .B(stable_counting), .C(stable_counting_N_2131), 
         .Z(n14472)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16415_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_186 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4_adj_2425)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_186.init = 16'h7bde;
    LUT4 i2407_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2407_2_lut.init = 16'h6666;
    LUT4 i2409_2_lut_rep_381 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21482)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2409_2_lut_rep_381.init = 16'h8888;
    LUT4 i2414_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2414_2_lut_3_lut.init = 16'h7878;
    LUT4 i2416_2_lut_rep_356_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21457)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2416_2_lut_rep_356_3_lut.init = 16'h8080;
    LUT4 i2423_2_lut_rep_338_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21439)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2423_2_lut_rep_338_3_lut_4_lut.init = 16'h8000;
    LUT4 i2421_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2421_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21414), .SP(stable_counting), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21423), .SP(stable_counting), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX stable_count__i0 (.D(n63[0]), .SP(stable_counting), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22206), .SP(clk_1mhz_enable_185), .CD(n14472), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    LUT4 i2435_2_lut_rep_313_3_lut_4_lut (.A(stable_count[3]), .B(n21457), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21414)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2435_2_lut_rep_313_3_lut_4_lut.init = 16'h78f0;
    
endmodule
//
// Verilog Description of module COMMUTATION_U6
//

module COMMUTATION_U6 (MB_m3_c_0, clkout_c, MC_m3_c_0, n21485, dir_m3, 
            hallsense_m3, LED3_c, enable_m3, PWM_m3, MA_m3_c_1, n21452, 
            MA_m3_c_0, n14203, MC_m3_c_1, n3139, MB_m3_c_1, n3105);
    output MB_m3_c_0;
    input clkout_c;
    output MC_m3_c_0;
    output n21485;
    input dir_m3;
    input [2:0]hallsense_m3;
    input LED3_c;
    input enable_m3;
    input PWM_m3;
    output MA_m3_c_1;
    input n21452;
    output MA_m3_c_0;
    input n14203;
    output MC_m3_c_1;
    input n3139;
    output MB_m3_c_1;
    input n3105;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire [1:0]MospairB_1__N_2141;
    wire [1:0]MospairC_1__N_2143;
    
    wire n21501, n15951, n21163, n8;
    
    FD1S3AX MospairB_i1 (.D(MospairB_1__N_2141[0]), .CK(clkout_c), .Q(MB_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=345, LSE_RLINE=345 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3AX MospairC_i1 (.D(MospairC_1__N_2143[0]), .CK(clkout_c), .Q(MC_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=345, LSE_RLINE=345 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i1.GSR = "DISABLED";
    LUT4 n21485_bdd_4_lut (.A(n21485), .B(dir_m3), .C(hallsense_m3[2]), 
         .D(hallsense_m3[0]), .Z(n21501)) /* synthesis lut_function=(!((B ((D)+!C)+!B (C+!(D)))+!A)) */ ;
    defparam n21485_bdd_4_lut.init = 16'h0280;
    LUT4 i17239_2_lut_3_lut (.A(LED3_c), .B(enable_m3), .C(PWM_m3), .Z(n15951)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17239_2_lut_3_lut.init = 16'h0404;
    LUT4 gnd_bdd_2_lut_17318_3_lut (.A(LED3_c), .B(enable_m3), .C(n21163), 
         .Z(MospairB_1__N_2141[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam gnd_bdd_2_lut_17318_3_lut.init = 16'h4040;
    LUT4 i21_4_lut (.A(hallsense_m3[0]), .B(n21485), .C(hallsense_m3[1]), 
         .D(dir_m3), .Z(n8)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i21_4_lut.init = 16'h400a;
    FD1S3IX MospairA_i2 (.D(n21501), .CK(clkout_c), .CD(n21452), .Q(MA_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=345, LSE_RLINE=345 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i2.GSR = "DISABLED";
    LUT4 PWM_m3_bdd_4_lut (.A(PWM_m3), .B(hallsense_m3[1]), .C(hallsense_m3[2]), 
         .D(dir_m3), .Z(n21163)) /* synthesis lut_function=((B (C+(D))+!B !(C (D)))+!A) */ ;
    defparam PWM_m3_bdd_4_lut.init = 16'hdff7;
    FD1S3JX MospairA_i1 (.D(n15951), .CK(clkout_c), .PD(n14203), .Q(MA_m3_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=345, LSE_RLINE=345 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i1.GSR = "DISABLED";
    FD1S3IX MospairC_i2 (.D(n21485), .CK(clkout_c), .CD(n3139), .Q(MC_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=345, LSE_RLINE=345 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n21485), .CK(clkout_c), .CD(n3105), .Q(MB_m3_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=345, LSE_RLINE=345 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i17170_2_lut_rep_384 (.A(LED3_c), .B(enable_m3), .Z(n21485)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17170_2_lut_rep_384.init = 16'h4444;
    LUT4 i17226_3_lut_4_lut (.A(LED3_c), .B(enable_m3), .C(n8), .D(PWM_m3), 
         .Z(MospairC_1__N_2143[0])) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17226_3_lut_4_lut.init = 16'h0444;
    
endmodule
//
// Verilog Description of module HALL_U3
//

module HALL_U3 (clk_1mhz, \speed_m3[0] , hallsense_m3, clkout_c_enable_362, 
            H_A_m3_c, H_B_m3_c, H_C_m3_c, \speed_m3[1] , \speed_m3[2] , 
            \speed_m3[3] , \speed_m3[4] , \speed_m3[5] , \speed_m3[6] , 
            \speed_m3[7] , \speed_m3[8] , \speed_m3[9] , \speed_m3[10] , 
            \speed_m3[11] , \speed_m3[12] , \speed_m3[13] , \speed_m3[14] , 
            \speed_m3[15] , \speed_m3[16] , \speed_m3[17] , \speed_m3[18] , 
            \speed_m3[19] , GND_net, n22206);
    input clk_1mhz;
    output \speed_m3[0] ;
    output [2:0]hallsense_m3;
    input clkout_c_enable_362;
    input H_A_m3_c;
    input H_B_m3_c;
    input H_C_m3_c;
    output \speed_m3[1] ;
    output \speed_m3[2] ;
    output \speed_m3[3] ;
    output \speed_m3[4] ;
    output \speed_m3[5] ;
    output \speed_m3[6] ;
    output \speed_m3[7] ;
    output \speed_m3[8] ;
    output \speed_m3[9] ;
    output \speed_m3[10] ;
    output \speed_m3[11] ;
    output \speed_m3[12] ;
    output \speed_m3[13] ;
    output \speed_m3[14] ;
    output \speed_m3[15] ;
    output \speed_m3[16] ;
    output \speed_m3[17] ;
    output \speed_m3[18] ;
    output \speed_m3[19] ;
    input GND_net;
    input n22206;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire stable_counting, n14454, n21483;
    wire [19:0]speedt_19__N_2049;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4626;
    wire [19:0]count_19__N_2069;
    
    wire hall3_lat;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_183, n18860, n19787, hall3_old, clk_1mhz_enable_184, 
        n19, n19588, n24, n20, hall1_old, hall2_old, hall1_lat, 
        hall2_lat, n22, n16, n11572, n11570, n19829, n19913, n19827, 
        n19895, n19835;
    wire [6:0]n63;
    
    wire n19577, n19654, n12, stable_counting_N_2131, n21415, n21479, 
        n21459, n4, n4_adj_2424, n21435, n21455, n18313, n18312, 
        n18311, n18310, n18309, n18308, n18307, n18306, n18305, 
        n18304;
    
    FD1P3IX stable_count__i0 (.D(n21483), .SP(stable_counting), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_2049[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_19__N_2069[0]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2069[0]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    LUT4 i17257_4_lut (.A(n18860), .B(n19787), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_184)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17257_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut (.A(n19), .B(n19588), .C(n24), .D(n20), .Z(n18860)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i16336_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19787)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16336_4_lut.init = 16'h7bde;
    LUT4 i6_2_lut (.A(count[17]), .B(count[12]), .Z(n19)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i11_4_lut (.A(count[5]), .B(n22), .C(n16), .D(count[16]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut (.A(count[14]), .B(count[19]), .C(count[11]), .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i7_3_lut.init = 16'hfefe;
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    LUT4 i9_4_lut (.A(count[15]), .B(count[18]), .C(count[1]), .D(count[4]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i9_4_lut.init = 16'hfffe;
    FD1P3AX hall1_lat_57 (.D(H_A_m3_c), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    FD1P3AX hall2_lat_58 (.D(H_B_m3_c), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m3_c), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    LUT4 i3_2_lut (.A(count[6]), .B(count[7]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(87[7:19])
    defparam i3_2_lut.init = 16'heeee;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2049[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2049[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2049[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2049[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2049[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2049[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2049[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2049[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2049[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2049[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2049[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2049[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2049[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2049[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2049[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2049[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2049[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2049[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2049[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11572), .B(n11570), .C(count_19__N_2069[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2049[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_179 (.A(n19588), .B(n19829), .C(n19913), .D(n19827), 
         .Z(n11572)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_179.init = 16'h0002;
    LUT4 i16377_2_lut (.A(count[18]), .B(count[1]), .Z(n19829)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16377_2_lut.init = 16'heeee;
    LUT4 i16461_4_lut (.A(count[7]), .B(n19895), .C(n19835), .D(count[15]), 
         .Z(n19913)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16461_4_lut.init = 16'hfffe;
    LUT4 i16375_3_lut (.A(count[5]), .B(count[17]), .C(count[16]), .Z(n19827)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i16375_3_lut.init = 16'hfefe;
    LUT4 i16443_4_lut (.A(count[11]), .B(count[12]), .C(count[4]), .D(count[6]), 
         .Z(n19895)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16443_4_lut.init = 16'hfffe;
    LUT4 i16383_2_lut (.A(count[19]), .B(count[14]), .Z(n19835)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16383_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(n63[4]), .B(stable_count[0]), .C(n19577), .D(n19654), 
         .Z(n11570)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i6_4_lut (.A(count[10]), .B(n12), .C(count[9]), .D(count[2]), 
         .Z(n19588)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[3]), .B(count[8]), .C(count[13]), .D(count[0]), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i2295_2_lut (.A(stable_counting), .B(stable_counting_N_2131), .Z(n4626)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2295_2_lut.init = 16'h8888;
    FD1P3AX speed__i2 (.D(speedt_19__N_2049[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2049[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2049[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2049[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2049[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2049[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2049[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2049[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m3[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2049[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2049[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2049[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2049[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2049[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2049[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2049[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2049[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2049[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2049[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2049[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m3[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(count_19__N_2069[1]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2069[2]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2069[3]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2069[4]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2069[5]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2069[6]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2069[7]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2069[8]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2069[9]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2069[10]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2069[11]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2069[12]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2069[13]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2069[14]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2069[15]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2069[16]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2069[17]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2069[18]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2069[19]), .CK(clk_1mhz), .CD(n4626), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n63[6]), .B(n63[3]), .C(n21415), .D(n63[2]), 
         .Z(n19577)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2069[1]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2069[2]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2069[3]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2069[4]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2069[5]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2069[6]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2069[7]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2069[8]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2069[9]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2069[10]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2069[11]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2069[12]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2069[13]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2069[14]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2069[15]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2069[16]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2069[17]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2069[18]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2069[19]), .SP(clk_1mhz_enable_183), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    LUT4 i2528_2_lut_3_lut_4_lut (.A(stable_count[2]), .B(n21479), .C(stable_count[4]), 
         .D(stable_count[3]), .Z(n63[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2528_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i16411_3_lut (.A(n21459), .B(stable_counting), .C(stable_counting_N_2131), 
         .Z(n14454)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16411_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_180 (.A(hall2_old), .B(hall1_old), .C(hall2_lat), 
         .D(hall1_lat), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_180.init = 16'h7bde;
    LUT4 i1_4_lut_adj_181 (.A(n63[2]), .B(n19654), .C(n63[4]), .D(n4_adj_2424), 
         .Z(stable_counting_N_2131)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_181.init = 16'h0004;
    LUT4 i11561_4_lut (.A(n11572), .B(n11570), .C(stable_counting), .D(stable_counting_N_2131), 
         .Z(clk_1mhz_enable_183)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11561_4_lut.init = 16'hcaea;
    LUT4 i2507_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2507_2_lut.init = 16'h6666;
    LUT4 i2542_3_lut_4_lut (.A(stable_count[4]), .B(n21435), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2542_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2_3_lut_rep_358 (.A(hall3_old), .B(n4), .C(hall3_lat), .Z(n21459)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_358.init = 16'hdede;
    LUT4 i1_2_lut_4_lut_adj_182 (.A(hall3_old), .B(n4), .C(hall3_lat), 
         .D(n63[1]), .Z(n19654)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_182.init = 16'h2100;
    LUT4 i2509_2_lut_rep_378 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21479)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2509_2_lut_rep_378.init = 16'h8888;
    LUT4 i2514_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2514_2_lut_3_lut.init = 16'h7878;
    LUT4 i2516_2_lut_rep_354_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21455)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2516_2_lut_rep_354_3_lut.init = 16'h8080;
    LUT4 i2523_2_lut_rep_334_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21435)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2523_2_lut_rep_334_3_lut_4_lut.init = 16'h8000;
    LUT4 i2521_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2521_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18313), 
          .S0(count_19__N_2069[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18312), .COUT(n18313), .S0(count_19__N_2069[17]), .S1(count_19__N_2069[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18311), .COUT(n18312), .S0(count_19__N_2069[15]), .S1(count_19__N_2069[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18310), .COUT(n18311), .S0(count_19__N_2069[13]), .S1(count_19__N_2069[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18309), .COUT(n18310), .S0(count_19__N_2069[11]), .S1(count_19__N_2069[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18308), .COUT(n18309), .S0(count_19__N_2069[9]), .S1(count_19__N_2069[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18307), 
          .COUT(n18308), .S0(count_19__N_2069[7]), .S1(count_19__N_2069[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18306), 
          .COUT(n18307), .S0(count_19__N_2069[5]), .S1(count_19__N_2069[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    LUT4 i2535_2_lut_rep_314_3_lut_4_lut (.A(stable_count[3]), .B(n21455), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21415)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2535_2_lut_rep_314_3_lut_4_lut.init = 16'h78f0;
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18305), 
          .COUT(n18306), .S0(count_19__N_2069[3]), .S1(count_19__N_2069[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18304), 
          .COUT(n18305), .S0(count_19__N_2069[1]), .S1(count_19__N_2069[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18304), 
          .S1(count_19__N_2069[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    LUT4 i2505_1_lut_rep_382 (.A(stable_count[0]), .Z(n21483)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2505_1_lut_rep_382.init = 16'h5555;
    LUT4 i1_2_lut_4_lut_4_lut (.A(stable_count[0]), .B(n21415), .C(n63[3]), 
         .D(n63[6]), .Z(n4_adj_2424)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_4_lut_4_lut.init = 16'hfffd;
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21415), .SP(stable_counting), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n63[4]), .SP(stable_counting), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22206), .SP(clk_1mhz_enable_184), .CD(n14454), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=342, LSE_RLINE=342 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module COMMUTATION
//

module COMMUTATION (MB_m4_c_0, clkout_c, MC_m4_c_0, n21484, dir_m4, 
            hallsense_m4, PWM_m4, MA_m4_c_1, n21449, LED4_c, enable_m4, 
            MC_m4_c_1, n3241, MB_m4_c_1, n3207, MA_m4_c_0, n14208);
    output MB_m4_c_0;
    input clkout_c;
    output MC_m4_c_0;
    output n21484;
    input dir_m4;
    input [2:0]hallsense_m4;
    input PWM_m4;
    output MA_m4_c_1;
    input n21449;
    input LED4_c;
    input enable_m4;
    output MC_m4_c_1;
    input n3241;
    output MB_m4_c_1;
    input n3207;
    output MA_m4_c_0;
    input n14208;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    wire [1:0]MospairB_1__N_2141;
    wire [1:0]MospairC_1__N_2143;
    
    wire n21500, n21147, n8, n15947;
    
    FD1S3AX MospairB_i1 (.D(MospairB_1__N_2141[0]), .CK(clkout_c), .Q(MB_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i1.GSR = "DISABLED";
    FD1S3AX MospairC_i1 (.D(MospairC_1__N_2143[0]), .CK(clkout_c), .Q(MC_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i1.GSR = "DISABLED";
    LUT4 n21484_bdd_4_lut (.A(n21484), .B(dir_m4), .C(hallsense_m4[2]), 
         .D(hallsense_m4[0]), .Z(n21500)) /* synthesis lut_function=(!((B ((D)+!C)+!B (C+!(D)))+!A)) */ ;
    defparam n21484_bdd_4_lut.init = 16'h0280;
    LUT4 PWM_m4_bdd_4_lut (.A(PWM_m4), .B(hallsense_m4[1]), .C(hallsense_m4[2]), 
         .D(dir_m4), .Z(n21147)) /* synthesis lut_function=((B (C+(D))+!B !(C (D)))+!A) */ ;
    defparam PWM_m4_bdd_4_lut.init = 16'hdff7;
    LUT4 i21_4_lut (.A(hallsense_m4[0]), .B(n21484), .C(hallsense_m4[1]), 
         .D(dir_m4), .Z(n8)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i21_4_lut.init = 16'h400a;
    FD1S3IX MospairA_i2 (.D(n21500), .CK(clkout_c), .CD(n21449), .Q(MA_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i2.GSR = "DISABLED";
    LUT4 i17179_2_lut_rep_383 (.A(LED4_c), .B(enable_m4), .Z(n21484)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17179_2_lut_rep_383.init = 16'h4444;
    LUT4 i17222_3_lut_4_lut (.A(LED4_c), .B(enable_m4), .C(n8), .D(PWM_m4), 
         .Z(MospairC_1__N_2143[0])) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17222_3_lut_4_lut.init = 16'h0444;
    FD1S3IX MospairC_i2 (.D(n21484), .CK(clkout_c), .CD(n3241), .Q(MC_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairC_i2.GSR = "DISABLED";
    FD1S3IX MospairB_i2 (.D(n21484), .CK(clkout_c), .CD(n3207), .Q(MB_m4_c_1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairB_i2.GSR = "DISABLED";
    LUT4 i17237_2_lut_3_lut (.A(LED4_c), .B(enable_m4), .C(PWM_m4), .Z(n15947)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam i17237_2_lut_3_lut.init = 16'h0404;
    LUT4 gnd_bdd_2_lut_17317_3_lut (.A(LED4_c), .B(enable_m4), .C(n21147), 
         .Z(MospairB_1__N_2141[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(69[3] 188[10])
    defparam gnd_bdd_2_lut_17317_3_lut.init = 16'h4040;
    FD1S3JX MospairA_i1 (.D(n15947), .CK(clkout_c), .PD(n14208), .Q(MA_m4_c_0)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=24, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/commutation.vhd(67[2] 189[9])
    defparam MospairA_i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AVG_SPEED
//

module AVG_SPEED (\speed_avg_m4[0] , clk_1mhz, \speed_m4[0] , \speed_avg_m4[1] , 
            \speed_m4[1] , \speed_avg_m4[2] , \speed_m4[2] , \speed_avg_m4[3] , 
            \speed_m4[3] , \speed_avg_m4[4] , \speed_m4[4] , \speed_avg_m4[5] , 
            \speed_m4[5] , \speed_avg_m4[6] , \speed_m4[6] , \speed_avg_m4[7] , 
            \speed_m4[7] , \speed_avg_m4[8] , \speed_m4[8] , \speed_avg_m4[9] , 
            \speed_m4[9] , \speed_avg_m4[10] , \speed_m4[10] , \speed_avg_m4[11] , 
            \speed_m4[11] , \speed_avg_m4[12] , \speed_m4[12] , \speed_avg_m4[13] , 
            \speed_m4[13] , \speed_avg_m4[14] , \speed_m4[14] , \speed_avg_m4[15] , 
            \speed_m4[15] , \speed_avg_m4[16] , \speed_m4[16] , \speed_avg_m4[17] , 
            \speed_m4[17] , \speed_avg_m4[18] , \speed_m4[18] , \speed_avg_m4[19] , 
            \speed_m4[19] , GND_net);
    output \speed_avg_m4[0] ;
    input clk_1mhz;
    input \speed_m4[0] ;
    output \speed_avg_m4[1] ;
    input \speed_m4[1] ;
    output \speed_avg_m4[2] ;
    input \speed_m4[2] ;
    output \speed_avg_m4[3] ;
    input \speed_m4[3] ;
    output \speed_avg_m4[4] ;
    input \speed_m4[4] ;
    output \speed_avg_m4[5] ;
    input \speed_m4[5] ;
    output \speed_avg_m4[6] ;
    input \speed_m4[6] ;
    output \speed_avg_m4[7] ;
    input \speed_m4[7] ;
    output \speed_avg_m4[8] ;
    input \speed_m4[8] ;
    output \speed_avg_m4[9] ;
    input \speed_m4[9] ;
    output \speed_avg_m4[10] ;
    input \speed_m4[10] ;
    output \speed_avg_m4[11] ;
    input \speed_m4[11] ;
    output \speed_avg_m4[12] ;
    input \speed_m4[12] ;
    output \speed_avg_m4[13] ;
    input \speed_m4[13] ;
    output \speed_avg_m4[14] ;
    input \speed_m4[14] ;
    output \speed_avg_m4[15] ;
    input \speed_m4[15] ;
    output \speed_avg_m4[16] ;
    input \speed_m4[16] ;
    output \speed_avg_m4[17] ;
    input \speed_m4[17] ;
    output \speed_avg_m4[18] ;
    input \speed_m4[18] ;
    output \speed_avg_m4[19] ;
    input \speed_m4[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_164;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n19839, n6, n18373, n18372, n18371;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m4[0] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2138__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_164), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138__i0.GSR = "DISABLED";
    LUT4 i17242_4_lut (.A(clk_cnt[0]), .B(n19839), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_164)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17242_4_lut.init = 16'h0004;
    LUT4 i16387_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n19839)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16387_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m4[1] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m4[2] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m4[3] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m4[4] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m4[5] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m4[6] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m4[7] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m4[8] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m4[9] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m4[10] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m4[11] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m4[12] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m4[13] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m4[14] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m4[15] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m4[16] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m4[17] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m4[18] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m4[19] ), .SP(clk_1mhz_enable_164), 
            .CK(clk_1mhz), .Q(\speed_avg_m4[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=370, LSE_RLINE=370 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    CCU2D clk_cnt_2138_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18373), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2138_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2138_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2138_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2138_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18372), .COUT(n18373), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2138_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2138_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2138_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2138_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18371), .COUT(n18372), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2138_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2138_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2138_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2138_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18371), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2138_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2138_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2138_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2138__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_164), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2138__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_164), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2138__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_164), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2138__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_164), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2138__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_164), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2138__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_164), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2138__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module SPI
//

module SPI (GND_net, clkout_c, MISO_N_816, n22211, speed_set_m2, speed_set_m4, 
            speed_set_m1, enable_m1, enable_m2, enable_m3, enable_m4, 
            clkout_c_enable_362, CS_c, SCK_c, MOSI_c, clkout_c_enable_266, 
            rst, n5199, speed_set_m3);
    input GND_net;
    input clkout_c;
    output MISO_N_816;
    input n22211;
    output [20:0]speed_set_m2;
    output [20:0]speed_set_m4;
    output [20:0]speed_set_m1;
    output enable_m1;
    output enable_m2;
    output enable_m3;
    output enable_m4;
    input clkout_c_enable_362;
    input CS_c;
    input SCK_c;
    input MOSI_c;
    input clkout_c_enable_266;
    input rst;
    output n5199;
    output [20:0]speed_set_m3;
    
    wire clkout_c /* synthesis SET_AS_NETWORK=clkout_c, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(44[2:8])
    
    wire n18475;
    wire [95:0]recv_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(68[10:21])
    
    wire n18476, n18474, n18473, n18472;
    wire [95:0]temp_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(70[10:21])
    
    wire clkout_c_enable_348;
    wire [95:0]n193;
    
    wire MISO_N_862, SCKold, CSlatched, SCKlatched, clkout_c_enable_60, 
        n14258;
    wire [95:0]send_buffer;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(67[10:21])
    
    wire n21454, n21456;
    wire [95:0]send_buffer_95__N_442;
    
    wire n14218, n14278, enable_m1_N_825, enable_m1_N_819, enable_m2_N_827, 
        enable_m3_N_834, enable_m4_N_841, CSold, n22207, MISO_N_817, 
        n21481, n18515, n3372, MISOb, MISOb_N_852, clkout_c_enable_107, 
        n3396, n39, n40, n36, n28, n38, n32, n34, n24, n3492, 
        n3468, n39_adj_2392, n40_adj_2393, n36_adj_2394, n28_adj_2395, 
        n38_adj_2396, n32_adj_2397, n34_adj_2398, n24_adj_2399, n3348, 
        n3324, n39_adj_2400, n40_adj_2401, n36_adj_2402, n28_adj_2403, 
        n38_adj_2404, n32_adj_2405, n34_adj_2406, n24_adj_2407, n3444, 
        n3420, n39_adj_2408, n40_adj_2409, n36_adj_2410, n28_adj_2411, 
        n38_adj_2412, n32_adj_2413, n34_adj_2414, n24_adj_2415, n18514, 
        n18513, n18512, n21480;
    wire [95:0]MISOb_N_858;
    
    wire MISOb_N_853, MISOb_N_857, n21442, n22208, n18511, n18510, 
        n18509, n18508, n18507, n18506, n18505, n18504, n18503, 
        n5197, n18502, n18501, n18500, n18499, n18498, n18429, 
        n18428, n18427, n18426, n18425, n18424, n18423, n18422, 
        n14238, n18623, n18622, n18621, n18620, n18619, n18618, 
        n18479, n18617, n18616, n18615, n18614, n18603, n18602, 
        n18601, n18600, n18599, n18598, n18597, n18596, n18595, 
        n18594, n18570, n18569, n18568, n18567, n18566, n18565, 
        n18564, n18563, n18562, n18561, n18560, n18559, n18558, 
        n18557, n18556, n18555, n18554, n18553, n18478, n18477;
    
    CCU2D add_15143_10 (.A0(recv_buffer[46]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[47]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18475), .COUT(n18476));
    defparam add_15143_10.INIT0 = 16'h5555;
    defparam add_15143_10.INIT1 = 16'h5aaa;
    defparam add_15143_10.INJECT1_0 = "NO";
    defparam add_15143_10.INJECT1_1 = "NO";
    CCU2D add_15143_8 (.A0(recv_buffer[44]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[45]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18474), .COUT(n18475));
    defparam add_15143_8.INIT0 = 16'h5aaa;
    defparam add_15143_8.INIT1 = 16'h5aaa;
    defparam add_15143_8.INJECT1_0 = "NO";
    defparam add_15143_8.INJECT1_1 = "NO";
    CCU2D add_15143_6 (.A0(recv_buffer[42]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[43]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18473), .COUT(n18474));
    defparam add_15143_6.INIT0 = 16'h5555;
    defparam add_15143_6.INIT1 = 16'h5555;
    defparam add_15143_6.INJECT1_0 = "NO";
    defparam add_15143_6.INJECT1_1 = "NO";
    CCU2D add_15143_4 (.A0(recv_buffer[40]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[41]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18472), .COUT(n18473));
    defparam add_15143_4.INIT0 = 16'h5aaa;
    defparam add_15143_4.INIT1 = 16'h5555;
    defparam add_15143_4.INJECT1_0 = "NO";
    defparam add_15143_4.INJECT1_1 = "NO";
    CCU2D add_15143_2 (.A0(recv_buffer[38]), .B0(recv_buffer[37]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[39]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18472));
    defparam add_15143_2.INIT0 = 16'h7000;
    defparam add_15143_2.INIT1 = 16'h5aaa;
    defparam add_15143_2.INJECT1_0 = "NO";
    defparam add_15143_2.INJECT1_1 = "NO";
    FD1P3AX temp_buffer_i0_i0 (.D(n193[0]), .SP(clkout_c_enable_348), .CK(clkout_c), 
            .Q(temp_buffer[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i0.GSR = "DISABLED";
    FD1S3AX MISO_128 (.D(MISO_N_862), .CK(clkout_c), .Q(MISO_N_816)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISO_128.GSR = "DISABLED";
    LUT4 i3_4_lut_rep_409 (.A(SCKold), .B(n22211), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_60)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut_rep_409.init = 16'h0400;
    FD1P3IX speed_set_m2_i0_i0 (.D(recv_buffer[54]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i0.GSR = "DISABLED";
    LUT4 i13248_2_lut_4_lut (.A(send_buffer[95]), .B(temp_buffer[95]), .C(n21454), 
         .D(n21456), .Z(send_buffer_95__N_442[95])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[3] 138[10])
    defparam i13248_2_lut_4_lut.init = 16'h00ca;
    FD1P3IX speed_set_m4_i0_i16 (.D(recv_buffer[28]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i0 (.D(recv_buffer[75]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i0.GSR = "DISABLED";
    FD1P3AX enable_m1_112 (.D(enable_m1_N_819), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m1_112.GSR = "ENABLED";
    FD1P3AX enable_m2_113 (.D(enable_m2_N_827), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m2_113.GSR = "ENABLED";
    FD1P3AX enable_m3_114 (.D(enable_m3_N_834), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m3_114.GSR = "ENABLED";
    FD1P3AX enable_m4_115 (.D(enable_m4_N_841), .SP(enable_m1_N_825), .CK(clkout_c), 
            .Q(enable_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam enable_m4_115.GSR = "ENABLED";
    FD1P3AX CSold_116 (.D(n22207), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(CSold));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_116.GSR = "DISABLED";
    FD1P3AX SCKold_117 (.D(SCKlatched), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(SCKold));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKold_117.GSR = "DISABLED";
    FD1P3AX CSlatched_118 (.D(CS_c), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(CSlatched));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_118.GSR = "DISABLED";
    FD1P3AX i104_129 (.D(n21481), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(MISO_N_817));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i104_129.GSR = "DISABLED";
    FD1P3AX SCKlatched_119 (.D(SCK_c), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(SCKlatched));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam SCKlatched_119.GSR = "DISABLED";
    FD1P3AX recv_buffer_rep_5__i0 (.D(recv_buffer[1]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(n193[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer_rep_5__i0.GSR = "DISABLED";
    CCU2D add_15142_21 (.A0(recv_buffer[74]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18515), .S1(n3372));
    defparam add_15142_21.INIT0 = 16'h5555;
    defparam add_15142_21.INIT1 = 16'h0000;
    defparam add_15142_21.INJECT1_0 = "NO";
    defparam add_15142_21.INJECT1_1 = "NO";
    FD1P3AX MISOb_121 (.D(MISOb_N_852), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(MISOb));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam MISOb_121.GSR = "DISABLED";
    FD1P3AX recv_buffer__i95 (.D(MOSI_c), .SP(clkout_c_enable_60), .CK(clkout_c), 
            .Q(recv_buffer[95])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i95.GSR = "DISABLED";
    FD1P3AX recv_buffer__i94 (.D(recv_buffer[95]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[94])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i94.GSR = "DISABLED";
    FD1P3AX recv_buffer__i93 (.D(recv_buffer[94]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i93.GSR = "DISABLED";
    FD1P3AX recv_buffer__i92 (.D(recv_buffer[93]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i92.GSR = "DISABLED";
    FD1P3AX recv_buffer__i91 (.D(recv_buffer[92]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i91.GSR = "DISABLED";
    FD1P3AX recv_buffer__i90 (.D(recv_buffer[91]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i90.GSR = "DISABLED";
    FD1P3AX recv_buffer__i89 (.D(recv_buffer[90]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i89.GSR = "DISABLED";
    FD1P3AX recv_buffer__i88 (.D(recv_buffer[89]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i88.GSR = "DISABLED";
    FD1P3AX recv_buffer__i87 (.D(recv_buffer[88]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i87.GSR = "DISABLED";
    FD1P3AX recv_buffer__i86 (.D(recv_buffer[87]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i86.GSR = "DISABLED";
    FD1P3AX recv_buffer__i85 (.D(recv_buffer[86]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i85.GSR = "DISABLED";
    FD1P3AX recv_buffer__i84 (.D(recv_buffer[85]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i84.GSR = "DISABLED";
    FD1P3AX recv_buffer__i83 (.D(recv_buffer[84]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i83.GSR = "DISABLED";
    FD1P3AX recv_buffer__i82 (.D(recv_buffer[83]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i82.GSR = "DISABLED";
    FD1P3AX recv_buffer__i81 (.D(recv_buffer[82]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i81.GSR = "DISABLED";
    FD1P3AX recv_buffer__i80 (.D(recv_buffer[81]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i80.GSR = "DISABLED";
    FD1P3AX recv_buffer__i79 (.D(recv_buffer[80]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i79.GSR = "DISABLED";
    FD1P3AX recv_buffer__i78 (.D(recv_buffer[79]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i78.GSR = "DISABLED";
    FD1P3AX recv_buffer__i77 (.D(recv_buffer[78]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i77.GSR = "DISABLED";
    FD1P3AX recv_buffer__i76 (.D(recv_buffer[77]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i76.GSR = "DISABLED";
    FD1P3AX recv_buffer__i75 (.D(recv_buffer[76]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i75.GSR = "DISABLED";
    FD1P3AX recv_buffer__i74 (.D(recv_buffer[75]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i74.GSR = "DISABLED";
    FD1P3AX recv_buffer__i73 (.D(recv_buffer[74]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i73.GSR = "DISABLED";
    FD1P3AX recv_buffer__i72 (.D(recv_buffer[73]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i72.GSR = "DISABLED";
    FD1P3AX recv_buffer__i71 (.D(recv_buffer[72]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i71.GSR = "DISABLED";
    FD1P3AX recv_buffer__i70 (.D(recv_buffer[71]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i70.GSR = "DISABLED";
    FD1P3AX recv_buffer__i69 (.D(recv_buffer[70]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i69.GSR = "DISABLED";
    FD1P3AX recv_buffer__i68 (.D(recv_buffer[69]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i68.GSR = "DISABLED";
    FD1P3AX recv_buffer__i67 (.D(recv_buffer[68]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i67.GSR = "DISABLED";
    FD1P3AX recv_buffer__i66 (.D(recv_buffer[67]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i66.GSR = "DISABLED";
    FD1P3AX recv_buffer__i65 (.D(recv_buffer[66]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i65.GSR = "DISABLED";
    FD1P3AX recv_buffer__i64 (.D(recv_buffer[65]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i64.GSR = "DISABLED";
    FD1P3AX recv_buffer__i63 (.D(recv_buffer[64]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i63.GSR = "DISABLED";
    FD1P3AX recv_buffer__i62 (.D(recv_buffer[63]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i62.GSR = "DISABLED";
    FD1P3AX recv_buffer__i61 (.D(recv_buffer[62]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i61.GSR = "DISABLED";
    FD1P3AX recv_buffer__i60 (.D(recv_buffer[61]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i60.GSR = "DISABLED";
    FD1P3AX recv_buffer__i59 (.D(recv_buffer[60]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i59.GSR = "DISABLED";
    FD1P3AX recv_buffer__i58 (.D(recv_buffer[59]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i58.GSR = "DISABLED";
    FD1P3AX recv_buffer__i57 (.D(recv_buffer[58]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i57.GSR = "DISABLED";
    FD1P3AX recv_buffer__i56 (.D(recv_buffer[57]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i56.GSR = "DISABLED";
    FD1P3AX recv_buffer__i55 (.D(recv_buffer[56]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i55.GSR = "DISABLED";
    FD1P3AX recv_buffer__i54 (.D(recv_buffer[55]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i54.GSR = "DISABLED";
    FD1P3AX recv_buffer__i53 (.D(recv_buffer[54]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i53.GSR = "DISABLED";
    FD1P3AX recv_buffer__i52 (.D(recv_buffer[53]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i52.GSR = "DISABLED";
    FD1P3AX recv_buffer__i51 (.D(recv_buffer[52]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i51.GSR = "DISABLED";
    FD1P3AX recv_buffer__i50 (.D(recv_buffer[51]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i50.GSR = "DISABLED";
    FD1P3AX recv_buffer__i49 (.D(recv_buffer[50]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i49.GSR = "DISABLED";
    FD1P3AX recv_buffer__i48 (.D(recv_buffer[49]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i48.GSR = "DISABLED";
    FD1P3AX recv_buffer__i47 (.D(recv_buffer[48]), .SP(clkout_c_enable_60), 
            .CK(clkout_c), .Q(recv_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i47.GSR = "DISABLED";
    FD1P3AX recv_buffer__i46 (.D(recv_buffer[47]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i46.GSR = "DISABLED";
    FD1P3AX recv_buffer__i45 (.D(recv_buffer[46]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i45.GSR = "DISABLED";
    FD1P3AX recv_buffer__i44 (.D(recv_buffer[45]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i44.GSR = "DISABLED";
    FD1P3AX recv_buffer__i43 (.D(recv_buffer[44]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i43.GSR = "DISABLED";
    FD1P3AX recv_buffer__i42 (.D(recv_buffer[43]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i42.GSR = "DISABLED";
    FD1P3AX recv_buffer__i41 (.D(recv_buffer[42]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i41.GSR = "DISABLED";
    FD1P3AX recv_buffer__i40 (.D(recv_buffer[41]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i40.GSR = "DISABLED";
    FD1P3AX recv_buffer__i39 (.D(recv_buffer[40]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i39.GSR = "DISABLED";
    FD1P3AX recv_buffer__i38 (.D(recv_buffer[39]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i38.GSR = "DISABLED";
    FD1P3AX recv_buffer__i37 (.D(recv_buffer[38]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i37.GSR = "DISABLED";
    FD1P3AX recv_buffer__i36 (.D(recv_buffer[37]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i36.GSR = "DISABLED";
    FD1P3AX recv_buffer__i35 (.D(recv_buffer[36]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i35.GSR = "DISABLED";
    FD1P3AX recv_buffer__i34 (.D(recv_buffer[35]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i34.GSR = "DISABLED";
    FD1P3AX recv_buffer__i33 (.D(recv_buffer[34]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i33.GSR = "DISABLED";
    FD1P3AX recv_buffer__i32 (.D(recv_buffer[33]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i32.GSR = "DISABLED";
    FD1P3AX recv_buffer__i31 (.D(recv_buffer[32]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i31.GSR = "DISABLED";
    FD1P3AX recv_buffer__i30 (.D(recv_buffer[31]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i30.GSR = "DISABLED";
    FD1P3AX recv_buffer__i29 (.D(recv_buffer[30]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i29.GSR = "DISABLED";
    FD1P3AX recv_buffer__i28 (.D(recv_buffer[29]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i28.GSR = "DISABLED";
    FD1P3AX recv_buffer__i27 (.D(recv_buffer[28]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i27.GSR = "DISABLED";
    FD1P3AX recv_buffer__i26 (.D(recv_buffer[27]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i26.GSR = "DISABLED";
    FD1P3AX recv_buffer__i25 (.D(recv_buffer[26]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i25.GSR = "DISABLED";
    FD1P3AX recv_buffer__i24 (.D(recv_buffer[25]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i24.GSR = "DISABLED";
    FD1P3AX recv_buffer__i23 (.D(recv_buffer[24]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i23.GSR = "DISABLED";
    FD1P3AX recv_buffer__i22 (.D(recv_buffer[23]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i22.GSR = "DISABLED";
    FD1P3AX recv_buffer__i21 (.D(recv_buffer[22]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i21.GSR = "DISABLED";
    FD1P3AX recv_buffer__i20 (.D(recv_buffer[21]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i20.GSR = "DISABLED";
    FD1P3AX recv_buffer__i19 (.D(recv_buffer[20]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i19.GSR = "DISABLED";
    FD1P3AX recv_buffer__i18 (.D(recv_buffer[19]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i18.GSR = "DISABLED";
    FD1P3AX recv_buffer__i17 (.D(recv_buffer[18]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i17.GSR = "DISABLED";
    FD1P3AX recv_buffer__i16 (.D(recv_buffer[17]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i16.GSR = "DISABLED";
    FD1P3AX recv_buffer__i15 (.D(recv_buffer[16]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i15.GSR = "DISABLED";
    FD1P3AX recv_buffer__i14 (.D(recv_buffer[15]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i14.GSR = "DISABLED";
    FD1P3AX recv_buffer__i13 (.D(recv_buffer[14]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i13.GSR = "DISABLED";
    FD1P3AX recv_buffer__i12 (.D(recv_buffer[13]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i12.GSR = "DISABLED";
    FD1P3AX recv_buffer__i11 (.D(recv_buffer[12]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i11.GSR = "DISABLED";
    FD1P3AX recv_buffer__i10 (.D(recv_buffer[11]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i10.GSR = "DISABLED";
    FD1P3AX recv_buffer__i9 (.D(recv_buffer[10]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i9.GSR = "DISABLED";
    FD1P3AX recv_buffer__i8 (.D(recv_buffer[9]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i8.GSR = "DISABLED";
    FD1P3AX recv_buffer__i7 (.D(recv_buffer[8]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i7.GSR = "DISABLED";
    FD1P3AX recv_buffer__i6 (.D(recv_buffer[7]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i6.GSR = "DISABLED";
    FD1P3AX recv_buffer__i5 (.D(recv_buffer[6]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i5.GSR = "DISABLED";
    FD1P3AX recv_buffer__i4 (.D(recv_buffer[5]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i4.GSR = "DISABLED";
    FD1P3AX recv_buffer__i3 (.D(recv_buffer[4]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i3.GSR = "DISABLED";
    FD1P3AX recv_buffer__i2 (.D(recv_buffer[3]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i2.GSR = "DISABLED";
    FD1P3AX recv_buffer__i1 (.D(recv_buffer[2]), .SP(clkout_c_enable_107), 
            .CK(clkout_c), .Q(recv_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam recv_buffer__i1.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i95 (.D(recv_buffer[95]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[95])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i95.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i94 (.D(recv_buffer[94]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[94])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i94.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i93 (.D(recv_buffer[93]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i93.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i92 (.D(recv_buffer[92]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i92.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i91 (.D(recv_buffer[91]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i91.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i90 (.D(recv_buffer[90]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i90.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i89 (.D(recv_buffer[89]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i89.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i88 (.D(recv_buffer[88]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i88.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i87 (.D(recv_buffer[87]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i87.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i86 (.D(recv_buffer[86]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i86.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i85 (.D(recv_buffer[85]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i85.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i84 (.D(recv_buffer[84]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i84.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i83 (.D(recv_buffer[83]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i83.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i82 (.D(recv_buffer[82]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i82.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i81 (.D(recv_buffer[81]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i81.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i80 (.D(recv_buffer[80]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i80.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i79 (.D(recv_buffer[79]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i79.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i78 (.D(recv_buffer[78]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i78.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i77 (.D(recv_buffer[77]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i77.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i76 (.D(recv_buffer[76]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i76.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i75 (.D(recv_buffer[75]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i75.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i74 (.D(recv_buffer[74]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i74.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i73 (.D(recv_buffer[73]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i73.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i72 (.D(recv_buffer[72]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i72.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i71 (.D(recv_buffer[71]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i71.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i70 (.D(recv_buffer[70]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i70.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i69 (.D(recv_buffer[69]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i69.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i68 (.D(recv_buffer[68]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i68.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i67 (.D(recv_buffer[67]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i67.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i66 (.D(recv_buffer[66]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i66.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i65 (.D(recv_buffer[65]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i65.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i64 (.D(recv_buffer[64]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i64.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i63 (.D(recv_buffer[63]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i63.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i62 (.D(recv_buffer[62]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i62.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i61 (.D(recv_buffer[61]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i61.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i60 (.D(recv_buffer[60]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i60.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i59 (.D(recv_buffer[59]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i59.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i58 (.D(recv_buffer[58]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i58.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i57 (.D(recv_buffer[57]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i57.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i56 (.D(recv_buffer[56]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i56.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i55 (.D(recv_buffer[55]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i55.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i54 (.D(recv_buffer[54]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i54.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i53 (.D(recv_buffer[53]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i53.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i52 (.D(recv_buffer[52]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i52.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i51 (.D(recv_buffer[51]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i51.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i50 (.D(recv_buffer[50]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i50.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i49 (.D(recv_buffer[49]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i49.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i48 (.D(recv_buffer[48]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i48.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i47 (.D(recv_buffer[47]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i47.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i46 (.D(recv_buffer[46]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i46.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i45 (.D(recv_buffer[45]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i45.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i44 (.D(recv_buffer[44]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i44.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i43 (.D(recv_buffer[43]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i43.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i42 (.D(recv_buffer[42]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i42.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i41 (.D(recv_buffer[41]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i41.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i40 (.D(recv_buffer[40]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i40.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i39 (.D(recv_buffer[39]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i39.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i38 (.D(recv_buffer[38]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i38.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i37 (.D(recv_buffer[37]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i37.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i36 (.D(recv_buffer[36]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i36.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i35 (.D(recv_buffer[35]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i35.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i34 (.D(recv_buffer[34]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i34.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i33 (.D(recv_buffer[33]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i33.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i32 (.D(recv_buffer[32]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i32.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i31 (.D(recv_buffer[31]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i31.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i30 (.D(recv_buffer[30]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i30.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i29 (.D(recv_buffer[29]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i29.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i28 (.D(recv_buffer[28]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i28.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i27 (.D(recv_buffer[27]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i27.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i26 (.D(recv_buffer[26]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i26.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i25 (.D(recv_buffer[25]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i25.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i24 (.D(recv_buffer[24]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i24.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i23 (.D(recv_buffer[23]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i23.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i22 (.D(recv_buffer[22]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i22.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i21 (.D(recv_buffer[21]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i21.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i20 (.D(recv_buffer[20]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i20.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i19 (.D(recv_buffer[19]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i19.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i18 (.D(recv_buffer[18]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i18.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i17 (.D(recv_buffer[17]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i17.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i16 (.D(recv_buffer[16]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i16.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i15 (.D(recv_buffer[15]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i15.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i14 (.D(recv_buffer[14]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i14.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i13 (.D(recv_buffer[13]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i13.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i12 (.D(recv_buffer[12]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i12.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i11 (.D(recv_buffer[11]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i11.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i10 (.D(recv_buffer[10]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i10.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i9 (.D(recv_buffer[9]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i9.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i8 (.D(recv_buffer[8]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i8.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i7 (.D(recv_buffer[7]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i6 (.D(recv_buffer[6]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i5 (.D(recv_buffer[5]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i5.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i4 (.D(recv_buffer[4]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i4.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i3 (.D(recv_buffer[3]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i2 (.D(recv_buffer[2]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX temp_buffer_i0_i1 (.D(recv_buffer[1]), .SP(clkout_c_enable_348), 
            .CK(clkout_c), .Q(temp_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam temp_buffer_i0_i1.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(n3396), .B(n3372), .C(n39), .D(n40), .Z(enable_m2_N_827)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i18_4_lut (.A(recv_buffer[67]), .B(n36), .C(n28), .D(recv_buffer[66]), 
         .Z(n39)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(recv_buffer[69]), .B(n38), .C(n32), .D(recv_buffer[64]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(recv_buffer[54]), .B(recv_buffer[61]), .C(recv_buffer[71]), 
         .D(recv_buffer[65]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(recv_buffer[55]), .B(recv_buffer[56]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(recv_buffer[62]), .B(n34), .C(n24), .D(recv_buffer[70]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut (.A(recv_buffer[60]), .B(recv_buffer[57]), .C(recv_buffer[68]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i13_4_lut (.A(recv_buffer[74]), .B(recv_buffer[73]), .C(recv_buffer[63]), 
         .D(recv_buffer[58]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(recv_buffer[72]), .B(recv_buffer[59]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i2_4_lut_adj_152 (.A(n3492), .B(n3468), .C(n39_adj_2392), .D(n40_adj_2393), 
         .Z(enable_m4_N_841)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_152.init = 16'h8880;
    LUT4 i18_4_lut_adj_153 (.A(recv_buffer[25]), .B(n36_adj_2394), .C(n28_adj_2395), 
         .D(recv_buffer[24]), .Z(n39_adj_2392)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_153.init = 16'hfffe;
    LUT4 i19_4_lut_adj_154 (.A(recv_buffer[27]), .B(n38_adj_2396), .C(n32_adj_2397), 
         .D(recv_buffer[22]), .Z(n40_adj_2393)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_154.init = 16'hfffe;
    LUT4 i15_4_lut_adj_155 (.A(recv_buffer[12]), .B(recv_buffer[19]), .C(recv_buffer[29]), 
         .D(recv_buffer[23]), .Z(n36_adj_2394)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_155.init = 16'hfffe;
    LUT4 i7_2_lut_adj_156 (.A(recv_buffer[13]), .B(recv_buffer[14]), .Z(n28_adj_2395)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_156.init = 16'heeee;
    LUT4 i17_4_lut_adj_157 (.A(recv_buffer[20]), .B(n34_adj_2398), .C(n24_adj_2399), 
         .D(recv_buffer[28]), .Z(n38_adj_2396)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_157.init = 16'hfffe;
    LUT4 i11_3_lut_adj_158 (.A(recv_buffer[18]), .B(recv_buffer[15]), .C(recv_buffer[26]), 
         .Z(n32_adj_2397)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_158.init = 16'hfefe;
    LUT4 i13_4_lut_adj_159 (.A(recv_buffer[32]), .B(recv_buffer[31]), .C(recv_buffer[21]), 
         .D(recv_buffer[16]), .Z(n34_adj_2398)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_159.init = 16'hfffe;
    LUT4 i3_2_lut_adj_160 (.A(recv_buffer[30]), .B(recv_buffer[17]), .Z(n24_adj_2399)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_160.init = 16'heeee;
    FD1P3AX send_buffer_i0_i1 (.D(send_buffer_95__N_442[1]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i1.GSR = "DISABLED";
    LUT4 i2_4_lut_adj_161 (.A(n3348), .B(n3324), .C(n39_adj_2400), .D(n40_adj_2401), 
         .Z(enable_m1_N_819)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_161.init = 16'h8880;
    LUT4 i18_4_lut_adj_162 (.A(recv_buffer[88]), .B(n36_adj_2402), .C(n28_adj_2403), 
         .D(recv_buffer[87]), .Z(n39_adj_2400)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_162.init = 16'hfffe;
    FD1P3AX send_buffer_i0_i2 (.D(send_buffer_95__N_442[2]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i3 (.D(send_buffer_95__N_442[3]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i4 (.D(send_buffer_95__N_442[4]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i4.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i5 (.D(send_buffer_95__N_442[5]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i5.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i6 (.D(send_buffer_95__N_442[6]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i7 (.D(send_buffer_95__N_442[7]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i8 (.D(send_buffer_95__N_442[8]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i8.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i9 (.D(send_buffer_95__N_442[9]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i9.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i10 (.D(send_buffer_95__N_442[10]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i10.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i11 (.D(send_buffer_95__N_442[11]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i11.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i12 (.D(send_buffer_95__N_442[12]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i12.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i13 (.D(send_buffer_95__N_442[13]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i13.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i14 (.D(send_buffer_95__N_442[14]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i14.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i15 (.D(send_buffer_95__N_442[15]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i15.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i16 (.D(send_buffer_95__N_442[16]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i16.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i17 (.D(send_buffer_95__N_442[17]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i17.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i18 (.D(send_buffer_95__N_442[18]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i18.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i19 (.D(send_buffer_95__N_442[19]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i19.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i20 (.D(send_buffer_95__N_442[20]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i20.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i21 (.D(send_buffer_95__N_442[21]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i21.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i22 (.D(send_buffer_95__N_442[22]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i22.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i23 (.D(send_buffer_95__N_442[23]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i23.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i24 (.D(send_buffer_95__N_442[24]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i24.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i25 (.D(send_buffer_95__N_442[25]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i25.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i26 (.D(send_buffer_95__N_442[26]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i26.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i27 (.D(send_buffer_95__N_442[27]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i27.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i28 (.D(send_buffer_95__N_442[28]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i28.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i29 (.D(send_buffer_95__N_442[29]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[29])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i29.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i30 (.D(send_buffer_95__N_442[30]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[30])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i30.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i31 (.D(send_buffer_95__N_442[31]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[31])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i31.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i32 (.D(send_buffer_95__N_442[32]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[32])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i32.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i33 (.D(send_buffer_95__N_442[33]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[33])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i33.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i34 (.D(send_buffer_95__N_442[34]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[34])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i34.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i35 (.D(send_buffer_95__N_442[35]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[35])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i35.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i36 (.D(send_buffer_95__N_442[36]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[36])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i36.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i37 (.D(send_buffer_95__N_442[37]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[37])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i37.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i38 (.D(send_buffer_95__N_442[38]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[38])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i38.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i39 (.D(send_buffer_95__N_442[39]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[39])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i39.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i40 (.D(send_buffer_95__N_442[40]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[40])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i40.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i41 (.D(send_buffer_95__N_442[41]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[41])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i41.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i42 (.D(send_buffer_95__N_442[42]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[42])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i42.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i43 (.D(send_buffer_95__N_442[43]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[43])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i43.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i44 (.D(send_buffer_95__N_442[44]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[44])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i44.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i45 (.D(send_buffer_95__N_442[45]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[45])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i45.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i46 (.D(send_buffer_95__N_442[46]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[46])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i46.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i47 (.D(send_buffer_95__N_442[47]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[47])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i47.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i48 (.D(send_buffer_95__N_442[48]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[48])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i48.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i49 (.D(send_buffer_95__N_442[49]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[49])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i49.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i50 (.D(send_buffer_95__N_442[50]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[50])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i50.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i51 (.D(send_buffer_95__N_442[51]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[51])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i51.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i52 (.D(send_buffer_95__N_442[52]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[52])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i52.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i53 (.D(send_buffer_95__N_442[53]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[53])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i53.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i54 (.D(send_buffer_95__N_442[54]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[54])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i54.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i55 (.D(send_buffer_95__N_442[55]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[55])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i55.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i56 (.D(send_buffer_95__N_442[56]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[56])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i56.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i57 (.D(send_buffer_95__N_442[57]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[57])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i57.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i58 (.D(send_buffer_95__N_442[58]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[58])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i58.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i59 (.D(send_buffer_95__N_442[59]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[59])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i59.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i60 (.D(send_buffer_95__N_442[60]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[60])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i60.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i61 (.D(send_buffer_95__N_442[61]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[61])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i61.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i62 (.D(send_buffer_95__N_442[62]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[62])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i62.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i63 (.D(send_buffer_95__N_442[63]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[63])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i63.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i64 (.D(send_buffer_95__N_442[64]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[64])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i64.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i65 (.D(send_buffer_95__N_442[65]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[65])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i65.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i66 (.D(send_buffer_95__N_442[66]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[66])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i66.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i67 (.D(send_buffer_95__N_442[67]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[67])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i67.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i68 (.D(send_buffer_95__N_442[68]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[68])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i68.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i69 (.D(send_buffer_95__N_442[69]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[69])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i69.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i70 (.D(send_buffer_95__N_442[70]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[70])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i70.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i71 (.D(send_buffer_95__N_442[71]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[71])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i71.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i72 (.D(send_buffer_95__N_442[72]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[72])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i72.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i73 (.D(send_buffer_95__N_442[73]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[73])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i73.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i74 (.D(send_buffer_95__N_442[74]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[74])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i74.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i75 (.D(send_buffer_95__N_442[75]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[75])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i75.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i76 (.D(send_buffer_95__N_442[76]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[76])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i76.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i77 (.D(send_buffer_95__N_442[77]), .SP(clkout_c_enable_266), 
            .CK(clkout_c), .Q(send_buffer[77])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i77.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i78 (.D(send_buffer_95__N_442[78]), .SP(clkout_c_enable_362), 
            .CK(clkout_c), .Q(send_buffer[78])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i78.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i79 (.D(send_buffer_95__N_442[79]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[79])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i79.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i80 (.D(send_buffer_95__N_442[80]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[80])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i80.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i81 (.D(send_buffer_95__N_442[81]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[81])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i81.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i82 (.D(send_buffer_95__N_442[82]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[82])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i82.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i83 (.D(send_buffer_95__N_442[83]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[83])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i83.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i84 (.D(send_buffer_95__N_442[84]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[84])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i84.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i85 (.D(send_buffer_95__N_442[85]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[85])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i85.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i86 (.D(send_buffer_95__N_442[86]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[86])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i86.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i87 (.D(send_buffer_95__N_442[87]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[87])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i87.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i88 (.D(send_buffer_95__N_442[88]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[88])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i88.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i89 (.D(send_buffer_95__N_442[89]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[89])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i89.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i90 (.D(send_buffer_95__N_442[90]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[90])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i90.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i91 (.D(send_buffer_95__N_442[91]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[91])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i91.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i92 (.D(send_buffer_95__N_442[92]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[92])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i92.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i93 (.D(send_buffer_95__N_442[93]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[93])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i93.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i94 (.D(send_buffer_95__N_442[94]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[94])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i94.GSR = "DISABLED";
    FD1P3AX send_buffer_i0_i95 (.D(send_buffer_95__N_442[95]), .SP(rst), 
            .CK(clkout_c), .Q(send_buffer[95])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam send_buffer_i0_i95.GSR = "DISABLED";
    LUT4 i19_4_lut_adj_163 (.A(recv_buffer[90]), .B(n38_adj_2404), .C(n32_adj_2405), 
         .D(recv_buffer[85]), .Z(n40_adj_2401)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_163.init = 16'hfffe;
    LUT4 i15_4_lut_adj_164 (.A(recv_buffer[75]), .B(recv_buffer[82]), .C(recv_buffer[92]), 
         .D(recv_buffer[86]), .Z(n36_adj_2402)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_164.init = 16'hfffe;
    LUT4 i7_2_lut_adj_165 (.A(recv_buffer[76]), .B(recv_buffer[77]), .Z(n28_adj_2403)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_165.init = 16'heeee;
    LUT4 i17_4_lut_adj_166 (.A(recv_buffer[83]), .B(n34_adj_2406), .C(n24_adj_2407), 
         .D(recv_buffer[91]), .Z(n38_adj_2404)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_166.init = 16'hfffe;
    LUT4 i11_3_lut_adj_167 (.A(recv_buffer[81]), .B(recv_buffer[78]), .C(recv_buffer[89]), 
         .Z(n32_adj_2405)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_167.init = 16'hfefe;
    LUT4 i13_4_lut_adj_168 (.A(recv_buffer[95]), .B(recv_buffer[94]), .C(recv_buffer[84]), 
         .D(recv_buffer[79]), .Z(n34_adj_2406)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_168.init = 16'hfffe;
    LUT4 i3_2_lut_adj_169 (.A(recv_buffer[93]), .B(recv_buffer[80]), .Z(n24_adj_2407)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_169.init = 16'heeee;
    LUT4 CSold_I_0_136_2_lut (.A(CSold), .B(CSlatched), .Z(enable_m1_N_825)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam CSold_I_0_136_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_170 (.A(n3444), .B(n3420), .C(n39_adj_2408), .D(n40_adj_2409), 
         .Z(enable_m3_N_834)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_170.init = 16'h8880;
    LUT4 i18_4_lut_adj_171 (.A(recv_buffer[46]), .B(n36_adj_2410), .C(n28_adj_2411), 
         .D(recv_buffer[45]), .Z(n39_adj_2408)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_171.init = 16'hfffe;
    LUT4 i19_4_lut_adj_172 (.A(recv_buffer[48]), .B(n38_adj_2412), .C(n32_adj_2413), 
         .D(recv_buffer[43]), .Z(n40_adj_2409)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_172.init = 16'hfffe;
    LUT4 i15_4_lut_adj_173 (.A(recv_buffer[33]), .B(recv_buffer[40]), .C(recv_buffer[50]), 
         .D(recv_buffer[44]), .Z(n36_adj_2410)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_173.init = 16'hfffe;
    LUT4 i7_2_lut_adj_174 (.A(recv_buffer[34]), .B(recv_buffer[35]), .Z(n28_adj_2411)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_174.init = 16'heeee;
    LUT4 i17_4_lut_adj_175 (.A(recv_buffer[41]), .B(n34_adj_2414), .C(n24_adj_2415), 
         .D(recv_buffer[49]), .Z(n38_adj_2412)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_175.init = 16'hfffe;
    LUT4 i11_3_lut_adj_176 (.A(recv_buffer[39]), .B(recv_buffer[36]), .C(recv_buffer[47]), 
         .Z(n32_adj_2413)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_176.init = 16'hfefe;
    LUT4 i13_4_lut_adj_177 (.A(recv_buffer[53]), .B(recv_buffer[52]), .C(recv_buffer[42]), 
         .D(recv_buffer[37]), .Z(n34_adj_2414)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_177.init = 16'hfffe;
    LUT4 i3_2_lut_adj_178 (.A(recv_buffer[51]), .B(recv_buffer[38]), .Z(n24_adj_2415)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_178.init = 16'heeee;
    LUT4 i3_4_lut (.A(SCKold), .B(n22211), .C(CSlatched), .D(SCKlatched), 
         .Z(clkout_c_enable_107)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam i3_4_lut.init = 16'h0400;
    CCU2D add_15142_19 (.A0(recv_buffer[72]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[73]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18514), .COUT(n18515));
    defparam add_15142_19.INIT0 = 16'hf555;
    defparam add_15142_19.INIT1 = 16'hf555;
    defparam add_15142_19.INJECT1_0 = "NO";
    defparam add_15142_19.INJECT1_1 = "NO";
    CCU2D add_15142_17 (.A0(recv_buffer[70]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[71]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18513), .COUT(n18514));
    defparam add_15142_17.INIT0 = 16'hf555;
    defparam add_15142_17.INIT1 = 16'hf555;
    defparam add_15142_17.INJECT1_0 = "NO";
    defparam add_15142_17.INJECT1_1 = "NO";
    CCU2D add_15142_15 (.A0(recv_buffer[68]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[69]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18512), .COUT(n18513));
    defparam add_15142_15.INIT0 = 16'hf555;
    defparam add_15142_15.INIT1 = 16'hf555;
    defparam add_15142_15.INJECT1_0 = "NO";
    defparam add_15142_15.INJECT1_1 = "NO";
    LUT4 SCKold_I_0_2_lut_rep_379 (.A(SCKold), .B(SCKlatched), .Z(n21480)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(193[8:45])
    defparam SCKold_I_0_2_lut_rep_379.init = 16'h2222;
    LUT4 MISOb_N_853_I_0_3_lut_4_lut (.A(SCKold), .B(SCKlatched), .C(MISOb_N_858[1]), 
         .D(MISOb_N_853), .Z(MISOb_N_857)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(193[8:45])
    defparam MISOb_N_853_I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 CSlatched_I_0_1_lut_rep_380 (.A(CSlatched), .Z(n21481)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam CSlatched_I_0_1_lut_rep_380.init = 16'h5555;
    LUT4 mux_9_i96_3_lut_rep_341_4_lut_4_lut (.A(n22207), .B(send_buffer[95]), 
         .C(temp_buffer[95]), .D(CSold), .Z(n21442)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i96_3_lut_rep_341_4_lut_4_lut.init = 16'hd8cc;
    LUT4 CSold_I_0_2_lut_rep_353_2_lut (.A(n22207), .B(n22208), .Z(n21454)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam CSold_I_0_2_lut_rep_353_2_lut.init = 16'h4444;
    LUT4 MISOb_I_0_3_lut_4_lut_4_lut (.A(n22207), .B(MISOb), .C(temp_buffer[0]), 
         .D(n22208), .Z(MISOb_N_853)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam MISOb_I_0_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i92_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[91]), .C(temp_buffer[91]), 
         .D(n22208), .Z(MISOb_N_858[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i2_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[1]), .C(temp_buffer[1]), 
         .D(n22208), .Z(MISOb_N_858[1])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i2_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i3_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[2]), .C(temp_buffer[2]), 
         .D(n22208), .Z(MISOb_N_858[2])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i3_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i93_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[92]), .C(temp_buffer[92]), 
         .D(n22208), .Z(MISOb_N_858[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i94_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[93]), .C(temp_buffer[93]), 
         .D(n22208), .Z(MISOb_N_858[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i95_3_lut_4_lut_4_lut (.A(CSlatched), .B(send_buffer[94]), 
         .C(temp_buffer[94]), .D(n22208), .Z(MISOb_N_858[94])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i95_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15142_13 (.A0(recv_buffer[66]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[67]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18511), .COUT(n18512));
    defparam add_15142_13.INIT0 = 16'hf555;
    defparam add_15142_13.INIT1 = 16'h0aaa;
    defparam add_15142_13.INJECT1_0 = "NO";
    defparam add_15142_13.INJECT1_1 = "NO";
    CCU2D add_15142_11 (.A0(recv_buffer[64]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[65]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18510), .COUT(n18511));
    defparam add_15142_11.INIT0 = 16'h0aaa;
    defparam add_15142_11.INIT1 = 16'hf555;
    defparam add_15142_11.INJECT1_0 = "NO";
    defparam add_15142_11.INJECT1_1 = "NO";
    LUT4 mux_9_i4_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[3]), .C(temp_buffer[3]), 
         .D(n22208), .Z(MISOb_N_858[3])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i4_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i5_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[4]), .C(temp_buffer[4]), 
         .D(n22208), .Z(MISOb_N_858[4])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i5_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i6_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[5]), .C(temp_buffer[5]), 
         .D(n22208), .Z(MISOb_N_858[5])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i6_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i7_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[6]), .C(temp_buffer[6]), 
         .D(n22208), .Z(MISOb_N_858[6])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i7_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i8_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[7]), .C(temp_buffer[7]), 
         .D(n22208), .Z(MISOb_N_858[7])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i8_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15142_9 (.A0(recv_buffer[62]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[63]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18509), .COUT(n18510));
    defparam add_15142_9.INIT0 = 16'h0aaa;
    defparam add_15142_9.INIT1 = 16'h0aaa;
    defparam add_15142_9.INJECT1_0 = "NO";
    defparam add_15142_9.INJECT1_1 = "NO";
    CCU2D add_15142_7 (.A0(recv_buffer[60]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[61]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18508), .COUT(n18509));
    defparam add_15142_7.INIT0 = 16'hf555;
    defparam add_15142_7.INIT1 = 16'hf555;
    defparam add_15142_7.INJECT1_0 = "NO";
    defparam add_15142_7.INJECT1_1 = "NO";
    LUT4 mux_9_i9_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[8]), .C(temp_buffer[8]), 
         .D(n22208), .Z(MISOb_N_858[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i10_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[9]), .C(temp_buffer[9]), 
         .D(n22208), .Z(MISOb_N_858[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i11_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[10]), .C(temp_buffer[10]), 
         .D(n22208), .Z(MISOb_N_858[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i12_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[11]), .C(temp_buffer[11]), 
         .D(n22208), .Z(MISOb_N_858[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i13_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[12]), .C(temp_buffer[12]), 
         .D(n22208), .Z(MISOb_N_858[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i14_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[13]), .C(temp_buffer[13]), 
         .D(n22208), .Z(MISOb_N_858[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i15_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[14]), .C(temp_buffer[14]), 
         .D(n22208), .Z(MISOb_N_858[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i16_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[15]), .C(temp_buffer[15]), 
         .D(n22208), .Z(MISOb_N_858[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i17_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[16]), .C(temp_buffer[16]), 
         .D(n22208), .Z(MISOb_N_858[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i18_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[17]), .C(temp_buffer[17]), 
         .D(n22208), .Z(MISOb_N_858[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i19_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[18]), .C(temp_buffer[18]), 
         .D(n22208), .Z(MISOb_N_858[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i20_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[19]), .C(temp_buffer[19]), 
         .D(n22208), .Z(MISOb_N_858[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i21_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[20]), .C(temp_buffer[20]), 
         .D(n22208), .Z(MISOb_N_858[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i22_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[21]), .C(temp_buffer[21]), 
         .D(n22208), .Z(MISOb_N_858[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i23_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[22]), .C(temp_buffer[22]), 
         .D(n22208), .Z(MISOb_N_858[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i24_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[23]), .C(temp_buffer[23]), 
         .D(n22208), .Z(MISOb_N_858[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i25_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[24]), .C(temp_buffer[24]), 
         .D(n22208), .Z(MISOb_N_858[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i26_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[25]), .C(temp_buffer[25]), 
         .D(n22208), .Z(MISOb_N_858[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i27_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[26]), .C(temp_buffer[26]), 
         .D(n22208), .Z(MISOb_N_858[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i28_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[27]), .C(temp_buffer[27]), 
         .D(n22208), .Z(MISOb_N_858[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i29_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[28]), .C(temp_buffer[28]), 
         .D(n22208), .Z(MISOb_N_858[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i30_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[29]), .C(temp_buffer[29]), 
         .D(n22208), .Z(MISOb_N_858[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i31_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[30]), .C(temp_buffer[30]), 
         .D(n22208), .Z(MISOb_N_858[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i32_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[31]), .C(temp_buffer[31]), 
         .D(n22208), .Z(MISOb_N_858[31])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i32_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i33_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[32]), .C(temp_buffer[32]), 
         .D(n22208), .Z(MISOb_N_858[32])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i33_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i34_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[33]), .C(temp_buffer[33]), 
         .D(n22208), .Z(MISOb_N_858[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i35_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[34]), .C(temp_buffer[34]), 
         .D(n22208), .Z(MISOb_N_858[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i36_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[35]), .C(temp_buffer[35]), 
         .D(n22208), .Z(MISOb_N_858[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i37_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[36]), .C(temp_buffer[36]), 
         .D(n22208), .Z(MISOb_N_858[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i38_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[37]), .C(temp_buffer[37]), 
         .D(n22208), .Z(MISOb_N_858[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i39_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[38]), .C(temp_buffer[38]), 
         .D(n22208), .Z(MISOb_N_858[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i40_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[39]), .C(temp_buffer[39]), 
         .D(n22208), .Z(MISOb_N_858[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i41_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[40]), .C(temp_buffer[40]), 
         .D(n22208), .Z(MISOb_N_858[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i42_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[41]), .C(temp_buffer[41]), 
         .D(n22208), .Z(MISOb_N_858[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i43_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[42]), .C(temp_buffer[42]), 
         .D(n22208), .Z(MISOb_N_858[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i44_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[43]), .C(temp_buffer[43]), 
         .D(n22208), .Z(MISOb_N_858[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i45_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[44]), .C(temp_buffer[44]), 
         .D(n22208), .Z(MISOb_N_858[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15142_5 (.A0(recv_buffer[58]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[59]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18507), .COUT(n18508));
    defparam add_15142_5.INIT0 = 16'h0aaa;
    defparam add_15142_5.INIT1 = 16'hf555;
    defparam add_15142_5.INJECT1_0 = "NO";
    defparam add_15142_5.INJECT1_1 = "NO";
    CCU2D add_15142_3 (.A0(recv_buffer[56]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[57]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18506), .COUT(n18507));
    defparam add_15142_3.INIT0 = 16'hf555;
    defparam add_15142_3.INIT1 = 16'hf555;
    defparam add_15142_3.INJECT1_0 = "NO";
    defparam add_15142_3.INJECT1_1 = "NO";
    CCU2D add_15142_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[54]), .B1(recv_buffer[55]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18506));
    defparam add_15142_1.INIT0 = 16'hF000;
    defparam add_15142_1.INIT1 = 16'ha666;
    defparam add_15142_1.INJECT1_0 = "NO";
    defparam add_15142_1.INJECT1_1 = "NO";
    LUT4 mux_9_i46_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[45]), .C(temp_buffer[45]), 
         .D(n22208), .Z(MISOb_N_858[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i47_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[46]), .C(temp_buffer[46]), 
         .D(n22208), .Z(MISOb_N_858[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i48_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[47]), .C(temp_buffer[47]), 
         .D(n22208), .Z(MISOb_N_858[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i49_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[48]), .C(temp_buffer[48]), 
         .D(n22208), .Z(MISOb_N_858[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i50_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[49]), .C(temp_buffer[49]), 
         .D(n22208), .Z(MISOb_N_858[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i51_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[50]), .C(temp_buffer[50]), 
         .D(n22208), .Z(MISOb_N_858[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i52_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[51]), .C(temp_buffer[51]), 
         .D(n22208), .Z(MISOb_N_858[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i53_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[52]), .C(temp_buffer[52]), 
         .D(n22208), .Z(MISOb_N_858[52])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i53_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i54_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[53]), .C(temp_buffer[53]), 
         .D(n22208), .Z(MISOb_N_858[53])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i54_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i55_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[54]), .C(temp_buffer[54]), 
         .D(n22208), .Z(MISOb_N_858[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i56_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[55]), .C(temp_buffer[55]), 
         .D(n22208), .Z(MISOb_N_858[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i57_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[56]), .C(temp_buffer[56]), 
         .D(n22208), .Z(MISOb_N_858[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i58_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[57]), .C(temp_buffer[57]), 
         .D(n22208), .Z(MISOb_N_858[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i59_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[58]), .C(temp_buffer[58]), 
         .D(n22208), .Z(MISOb_N_858[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i60_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[59]), .C(temp_buffer[59]), 
         .D(n22208), .Z(MISOb_N_858[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i61_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[60]), .C(temp_buffer[60]), 
         .D(n22208), .Z(MISOb_N_858[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i62_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[61]), .C(temp_buffer[61]), 
         .D(n22208), .Z(MISOb_N_858[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i63_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[62]), .C(temp_buffer[62]), 
         .D(n22208), .Z(MISOb_N_858[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i64_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[63]), .C(temp_buffer[63]), 
         .D(n22208), .Z(MISOb_N_858[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i65_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[64]), .C(temp_buffer[64]), 
         .D(n22208), .Z(MISOb_N_858[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i66_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[65]), .C(temp_buffer[65]), 
         .D(n22208), .Z(MISOb_N_858[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i67_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[66]), .C(temp_buffer[66]), 
         .D(n22208), .Z(MISOb_N_858[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i68_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[67]), .C(temp_buffer[67]), 
         .D(n22208), .Z(MISOb_N_858[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15122_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18505), 
          .S0(n3348));
    defparam add_15122_cout.INIT0 = 16'h0000;
    defparam add_15122_cout.INIT1 = 16'h0000;
    defparam add_15122_cout.INJECT1_0 = "NO";
    defparam add_15122_cout.INJECT1_1 = "NO";
    CCU2D add_15122_16 (.A0(recv_buffer[94]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[95]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18504), .COUT(n18505));
    defparam add_15122_16.INIT0 = 16'h5aaa;
    defparam add_15122_16.INIT1 = 16'h0aaa;
    defparam add_15122_16.INJECT1_0 = "NO";
    defparam add_15122_16.INJECT1_1 = "NO";
    LUT4 mux_9_i69_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[68]), .C(temp_buffer[68]), 
         .D(n22208), .Z(MISOb_N_858[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i70_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[69]), .C(temp_buffer[69]), 
         .D(n22208), .Z(MISOb_N_858[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i71_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[70]), .C(temp_buffer[70]), 
         .D(n22208), .Z(MISOb_N_858[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i72_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[71]), .C(temp_buffer[71]), 
         .D(n22208), .Z(MISOb_N_858[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i73_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[72]), .C(temp_buffer[72]), 
         .D(n22208), .Z(MISOb_N_858[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i74_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[73]), .C(temp_buffer[73]), 
         .D(n22208), .Z(MISOb_N_858[73])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i74_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i75_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[74]), .C(temp_buffer[74]), 
         .D(n22208), .Z(MISOb_N_858[74])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i75_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i76_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[75]), .C(temp_buffer[75]), 
         .D(n22208), .Z(MISOb_N_858[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i77_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[76]), .C(temp_buffer[76]), 
         .D(n22208), .Z(MISOb_N_858[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15122_14 (.A0(recv_buffer[92]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[93]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18503), .COUT(n18504));
    defparam add_15122_14.INIT0 = 16'h5aaa;
    defparam add_15122_14.INIT1 = 16'h5aaa;
    defparam add_15122_14.INJECT1_0 = "NO";
    defparam add_15122_14.INJECT1_1 = "NO";
    LUT4 mux_9_i78_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[77]), .C(temp_buffer[77]), 
         .D(n22208), .Z(MISOb_N_858[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i79_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[78]), .C(temp_buffer[78]), 
         .D(n22208), .Z(MISOb_N_858[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i80_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[79]), .C(temp_buffer[79]), 
         .D(n22208), .Z(MISOb_N_858[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i2764_2_lut (.A(MISO_N_816), .B(MISO_N_817), .Z(n5197)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    defparam i2764_2_lut.init = 16'h8888;
    LUT4 mux_9_i81_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[80]), .C(temp_buffer[80]), 
         .D(n22208), .Z(MISOb_N_858[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i82_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[81]), .C(temp_buffer[81]), 
         .D(n22208), .Z(MISOb_N_858[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i83_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[82]), .C(temp_buffer[82]), 
         .D(n22208), .Z(MISOb_N_858[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i84_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[83]), .C(temp_buffer[83]), 
         .D(n22208), .Z(MISOb_N_858[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i85_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[84]), .C(temp_buffer[84]), 
         .D(n22208), .Z(MISOb_N_858[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i86_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[85]), .C(temp_buffer[85]), 
         .D(n22208), .Z(MISOb_N_858[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i87_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[86]), .C(temp_buffer[86]), 
         .D(n22208), .Z(MISOb_N_858[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i88_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[87]), .C(temp_buffer[87]), 
         .D(n22208), .Z(MISOb_N_858[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i89_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[88]), .C(temp_buffer[88]), 
         .D(n22208), .Z(MISOb_N_858[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i90_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[89]), .C(temp_buffer[89]), 
         .D(n22208), .Z(MISOb_N_858[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_9_i91_3_lut_4_lut_4_lut (.A(n22207), .B(send_buffer[90]), .C(temp_buffer[90]), 
         .D(n22208), .Z(MISOb_N_858[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_9_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15122_12 (.A0(recv_buffer[90]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[91]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18502), .COUT(n18503));
    defparam add_15122_12.INIT0 = 16'h5aaa;
    defparam add_15122_12.INIT1 = 16'h5aaa;
    defparam add_15122_12.INJECT1_0 = "NO";
    defparam add_15122_12.INJECT1_1 = "NO";
    LUT4 i2976_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_853), .C(MISOb_N_858[1]), 
         .D(n21480), .Z(MISOb_N_852)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam i2976_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i2_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[1]), 
         .C(MISOb_N_858[2]), .D(n21480), .Z(send_buffer_95__N_442[1])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i2_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i3_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[2]), 
         .C(MISOb_N_858[3]), .D(n21480), .Z(send_buffer_95__N_442[2])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i3_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i4_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[3]), 
         .C(MISOb_N_858[4]), .D(n21480), .Z(send_buffer_95__N_442[3])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i4_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15122_10 (.A0(recv_buffer[88]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[89]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18501), .COUT(n18502));
    defparam add_15122_10.INIT0 = 16'h5555;
    defparam add_15122_10.INIT1 = 16'h5aaa;
    defparam add_15122_10.INJECT1_0 = "NO";
    defparam add_15122_10.INJECT1_1 = "NO";
    CCU2D add_15122_8 (.A0(recv_buffer[86]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[87]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18500), .COUT(n18501));
    defparam add_15122_8.INIT0 = 16'h5aaa;
    defparam add_15122_8.INIT1 = 16'h5aaa;
    defparam add_15122_8.INJECT1_0 = "NO";
    defparam add_15122_8.INJECT1_1 = "NO";
    LUT4 mux_52_i5_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[4]), 
         .C(MISOb_N_858[5]), .D(n21480), .Z(send_buffer_95__N_442[4])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i5_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i6_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[5]), 
         .C(MISOb_N_858[6]), .D(n21480), .Z(send_buffer_95__N_442[5])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i6_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i7_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[6]), 
         .C(MISOb_N_858[7]), .D(n21480), .Z(send_buffer_95__N_442[6])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i7_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i8_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[7]), 
         .C(MISOb_N_858[8]), .D(n21480), .Z(send_buffer_95__N_442[7])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i8_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15122_6 (.A0(recv_buffer[84]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[85]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18499), .COUT(n18500));
    defparam add_15122_6.INIT0 = 16'h5555;
    defparam add_15122_6.INIT1 = 16'h5555;
    defparam add_15122_6.INJECT1_0 = "NO";
    defparam add_15122_6.INJECT1_1 = "NO";
    LUT4 mux_52_i9_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[8]), 
         .C(MISOb_N_858[9]), .D(n21480), .Z(send_buffer_95__N_442[8])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i9_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i10_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[9]), 
         .C(MISOb_N_858[10]), .D(n21480), .Z(send_buffer_95__N_442[9])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i10_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i11_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[10]), 
         .C(MISOb_N_858[11]), .D(n21480), .Z(send_buffer_95__N_442[10])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i11_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i12_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[11]), 
         .C(MISOb_N_858[12]), .D(n21480), .Z(send_buffer_95__N_442[11])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i12_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i13_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[12]), 
         .C(MISOb_N_858[13]), .D(n21480), .Z(send_buffer_95__N_442[12])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i13_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i14_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[13]), 
         .C(MISOb_N_858[14]), .D(n21480), .Z(send_buffer_95__N_442[13])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i14_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15122_4 (.A0(recv_buffer[82]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[83]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18498), .COUT(n18499));
    defparam add_15122_4.INIT0 = 16'h5aaa;
    defparam add_15122_4.INIT1 = 16'h5555;
    defparam add_15122_4.INJECT1_0 = "NO";
    defparam add_15122_4.INJECT1_1 = "NO";
    CCU2D add_15122_2 (.A0(recv_buffer[80]), .B0(recv_buffer[79]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[81]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18498));
    defparam add_15122_2.INIT0 = 16'h7000;
    defparam add_15122_2.INIT1 = 16'h5aaa;
    defparam add_15122_2.INJECT1_0 = "NO";
    defparam add_15122_2.INJECT1_1 = "NO";
    LUT4 mux_52_i15_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[14]), 
         .C(MISOb_N_858[15]), .D(n21480), .Z(send_buffer_95__N_442[14])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i15_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i16_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[15]), 
         .C(MISOb_N_858[16]), .D(n21480), .Z(send_buffer_95__N_442[15])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i16_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i17_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[16]), 
         .C(MISOb_N_858[17]), .D(n21480), .Z(send_buffer_95__N_442[16])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i17_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i18_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[17]), 
         .C(MISOb_N_858[18]), .D(n21480), .Z(send_buffer_95__N_442[17])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i18_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i19_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[18]), 
         .C(MISOb_N_858[19]), .D(n21480), .Z(send_buffer_95__N_442[18])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i19_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i20_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[19]), 
         .C(MISOb_N_858[20]), .D(n21480), .Z(send_buffer_95__N_442[19])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i20_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i21_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[20]), 
         .C(MISOb_N_858[21]), .D(n21480), .Z(send_buffer_95__N_442[20])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i21_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i22_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[21]), 
         .C(MISOb_N_858[22]), .D(n21480), .Z(send_buffer_95__N_442[21])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i22_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i23_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[22]), 
         .C(MISOb_N_858[23]), .D(n21480), .Z(send_buffer_95__N_442[22])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i23_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i24_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[23]), 
         .C(MISOb_N_858[24]), .D(n21480), .Z(send_buffer_95__N_442[23])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i24_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i25_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[24]), 
         .C(MISOb_N_858[25]), .D(n21480), .Z(send_buffer_95__N_442[24])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i25_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i26_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[25]), 
         .C(MISOb_N_858[26]), .D(n21480), .Z(send_buffer_95__N_442[25])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i26_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i27_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[26]), 
         .C(MISOb_N_858[27]), .D(n21480), .Z(send_buffer_95__N_442[26])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i27_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i28_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[27]), 
         .C(MISOb_N_858[28]), .D(n21480), .Z(send_buffer_95__N_442[27])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i28_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i29_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[28]), 
         .C(MISOb_N_858[29]), .D(n21480), .Z(send_buffer_95__N_442[28])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i29_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i30_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[29]), 
         .C(MISOb_N_858[30]), .D(n21480), .Z(send_buffer_95__N_442[29])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i30_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i31_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[30]), 
         .C(MISOb_N_858[31]), .D(n21480), .Z(send_buffer_95__N_442[30])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i31_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i32_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[31]), 
         .C(MISOb_N_858[32]), .D(n21480), .Z(send_buffer_95__N_442[31])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i32_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i33_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[32]), 
         .C(MISOb_N_858[33]), .D(n21480), .Z(send_buffer_95__N_442[32])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i33_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i34_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[33]), 
         .C(MISOb_N_858[34]), .D(n21480), .Z(send_buffer_95__N_442[33])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i34_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i35_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[34]), 
         .C(MISOb_N_858[35]), .D(n21480), .Z(send_buffer_95__N_442[34])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i35_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i36_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[35]), 
         .C(MISOb_N_858[36]), .D(n21480), .Z(send_buffer_95__N_442[35])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i36_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i37_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[36]), 
         .C(MISOb_N_858[37]), .D(n21480), .Z(send_buffer_95__N_442[36])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i37_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i38_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[37]), 
         .C(MISOb_N_858[38]), .D(n21480), .Z(send_buffer_95__N_442[37])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i38_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i39_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[38]), 
         .C(MISOb_N_858[39]), .D(n21480), .Z(send_buffer_95__N_442[38])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i39_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i40_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[39]), 
         .C(MISOb_N_858[40]), .D(n21480), .Z(send_buffer_95__N_442[39])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i40_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i41_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[40]), 
         .C(MISOb_N_858[41]), .D(n21480), .Z(send_buffer_95__N_442[40])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i41_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i42_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[41]), 
         .C(MISOb_N_858[42]), .D(n21480), .Z(send_buffer_95__N_442[41])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i42_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i43_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[42]), 
         .C(MISOb_N_858[43]), .D(n21480), .Z(send_buffer_95__N_442[42])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i43_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i44_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[43]), 
         .C(MISOb_N_858[44]), .D(n21480), .Z(send_buffer_95__N_442[43])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i44_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i45_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[44]), 
         .C(MISOb_N_858[45]), .D(n21480), .Z(send_buffer_95__N_442[44])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i45_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i46_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[45]), 
         .C(MISOb_N_858[46]), .D(n21480), .Z(send_buffer_95__N_442[45])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i46_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i47_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[46]), 
         .C(MISOb_N_858[47]), .D(n21480), .Z(send_buffer_95__N_442[46])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i47_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i48_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[47]), 
         .C(MISOb_N_858[48]), .D(n21480), .Z(send_buffer_95__N_442[47])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i48_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i49_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[48]), 
         .C(MISOb_N_858[49]), .D(n21480), .Z(send_buffer_95__N_442[48])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i49_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i50_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[49]), 
         .C(MISOb_N_858[50]), .D(n21480), .Z(send_buffer_95__N_442[49])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i50_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i51_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[50]), 
         .C(MISOb_N_858[51]), .D(n21480), .Z(send_buffer_95__N_442[50])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i51_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i52_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[51]), 
         .C(MISOb_N_858[52]), .D(n21480), .Z(send_buffer_95__N_442[51])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i52_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i53_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[52]), 
         .C(MISOb_N_858[53]), .D(n21480), .Z(send_buffer_95__N_442[52])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i53_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i54_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[53]), 
         .C(MISOb_N_858[54]), .D(n21480), .Z(send_buffer_95__N_442[53])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i54_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i55_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[54]), 
         .C(MISOb_N_858[55]), .D(n21480), .Z(send_buffer_95__N_442[54])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i55_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i56_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[55]), 
         .C(MISOb_N_858[56]), .D(n21480), .Z(send_buffer_95__N_442[55])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i56_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i57_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[56]), 
         .C(MISOb_N_858[57]), .D(n21480), .Z(send_buffer_95__N_442[56])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i57_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i58_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[57]), 
         .C(MISOb_N_858[58]), .D(n21480), .Z(send_buffer_95__N_442[57])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i58_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i59_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[58]), 
         .C(MISOb_N_858[59]), .D(n21480), .Z(send_buffer_95__N_442[58])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i59_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i60_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[59]), 
         .C(MISOb_N_858[60]), .D(n21480), .Z(send_buffer_95__N_442[59])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i60_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i61_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[60]), 
         .C(MISOb_N_858[61]), .D(n21480), .Z(send_buffer_95__N_442[60])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i61_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i62_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[61]), 
         .C(MISOb_N_858[62]), .D(n21480), .Z(send_buffer_95__N_442[61])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i62_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i63_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[62]), 
         .C(MISOb_N_858[63]), .D(n21480), .Z(send_buffer_95__N_442[62])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i63_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i64_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[63]), 
         .C(MISOb_N_858[64]), .D(n21480), .Z(send_buffer_95__N_442[63])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i64_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i65_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[64]), 
         .C(MISOb_N_858[65]), .D(n21480), .Z(send_buffer_95__N_442[64])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i65_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i66_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[65]), 
         .C(MISOb_N_858[66]), .D(n21480), .Z(send_buffer_95__N_442[65])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i66_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i67_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[66]), 
         .C(MISOb_N_858[67]), .D(n21480), .Z(send_buffer_95__N_442[66])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i67_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i68_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[67]), 
         .C(MISOb_N_858[68]), .D(n21480), .Z(send_buffer_95__N_442[67])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i68_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i69_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[68]), 
         .C(MISOb_N_858[69]), .D(n21480), .Z(send_buffer_95__N_442[68])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i69_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i70_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[69]), 
         .C(MISOb_N_858[70]), .D(n21480), .Z(send_buffer_95__N_442[69])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i70_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i71_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[70]), 
         .C(MISOb_N_858[71]), .D(n21480), .Z(send_buffer_95__N_442[70])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i71_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i72_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[71]), 
         .C(MISOb_N_858[72]), .D(n21480), .Z(send_buffer_95__N_442[71])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i72_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i73_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[72]), 
         .C(MISOb_N_858[73]), .D(n21480), .Z(send_buffer_95__N_442[72])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i73_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i74_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[73]), 
         .C(MISOb_N_858[74]), .D(n21480), .Z(send_buffer_95__N_442[73])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i74_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i75_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[74]), 
         .C(MISOb_N_858[75]), .D(n21480), .Z(send_buffer_95__N_442[74])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i75_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i76_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[75]), 
         .C(MISOb_N_858[76]), .D(n21480), .Z(send_buffer_95__N_442[75])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i76_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i77_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[76]), 
         .C(MISOb_N_858[77]), .D(n21480), .Z(send_buffer_95__N_442[76])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i77_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i78_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[77]), 
         .C(MISOb_N_858[78]), .D(n21480), .Z(send_buffer_95__N_442[77])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i78_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i79_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[78]), 
         .C(MISOb_N_858[79]), .D(n21480), .Z(send_buffer_95__N_442[78])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i79_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i80_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[79]), 
         .C(MISOb_N_858[80]), .D(n21480), .Z(send_buffer_95__N_442[79])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i80_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i81_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[80]), 
         .C(MISOb_N_858[81]), .D(n21480), .Z(send_buffer_95__N_442[80])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i81_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i82_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[81]), 
         .C(MISOb_N_858[82]), .D(n21480), .Z(send_buffer_95__N_442[81])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i82_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i83_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[82]), 
         .C(MISOb_N_858[83]), .D(n21480), .Z(send_buffer_95__N_442[82])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i83_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i84_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[83]), 
         .C(MISOb_N_858[84]), .D(n21480), .Z(send_buffer_95__N_442[83])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i84_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i85_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[84]), 
         .C(MISOb_N_858[85]), .D(n21480), .Z(send_buffer_95__N_442[84])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i85_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i86_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[85]), 
         .C(MISOb_N_858[86]), .D(n21480), .Z(send_buffer_95__N_442[85])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i86_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i87_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[86]), 
         .C(MISOb_N_858[87]), .D(n21480), .Z(send_buffer_95__N_442[86])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i87_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i88_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[87]), 
         .C(MISOb_N_858[88]), .D(n21480), .Z(send_buffer_95__N_442[87])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i88_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i89_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[88]), 
         .C(MISOb_N_858[89]), .D(n21480), .Z(send_buffer_95__N_442[88])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i89_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i90_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[89]), 
         .C(MISOb_N_858[90]), .D(n21480), .Z(send_buffer_95__N_442[89])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i90_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i91_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[90]), 
         .C(MISOb_N_858[91]), .D(n21480), .Z(send_buffer_95__N_442[90])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i91_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D add_15136_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18429), 
          .S0(n3492));
    defparam add_15136_cout.INIT0 = 16'h0000;
    defparam add_15136_cout.INIT1 = 16'h0000;
    defparam add_15136_cout.INJECT1_0 = "NO";
    defparam add_15136_cout.INJECT1_1 = "NO";
    CCU2D add_15136_16 (.A0(recv_buffer[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[32]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18428), .COUT(n18429));
    defparam add_15136_16.INIT0 = 16'h5aaa;
    defparam add_15136_16.INIT1 = 16'h0aaa;
    defparam add_15136_16.INJECT1_0 = "NO";
    defparam add_15136_16.INJECT1_1 = "NO";
    LUT4 mux_52_i92_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[91]), 
         .C(MISOb_N_858[92]), .D(n21480), .Z(send_buffer_95__N_442[91])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i92_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i93_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[92]), 
         .C(MISOb_N_858[93]), .D(n21480), .Z(send_buffer_95__N_442[92])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i93_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i94_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[93]), 
         .C(MISOb_N_858[94]), .D(n21480), .Z(send_buffer_95__N_442[93])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i94_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 mux_52_i95_3_lut_4_lut_4_lut (.A(CSlatched), .B(MISOb_N_858[94]), 
         .C(n21442), .D(n21480), .Z(send_buffer_95__N_442[94])) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam mux_52_i95_3_lut_4_lut_4_lut.init = 16'hd8cc;
    LUT4 i163_2_lut_rep_355_3_lut_3_lut (.A(CSlatched), .B(SCKlatched), 
         .C(SCKold), .Z(n21456)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(117[26:41])
    defparam i163_2_lut_rep_355_3_lut_3_lut.init = 16'h1010;
    CCU2D add_15136_14 (.A0(recv_buffer[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18427), .COUT(n18428));
    defparam add_15136_14.INIT0 = 16'h5aaa;
    defparam add_15136_14.INIT1 = 16'h5aaa;
    defparam add_15136_14.INJECT1_0 = "NO";
    defparam add_15136_14.INJECT1_1 = "NO";
    CCU2D add_15136_12 (.A0(recv_buffer[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18426), .COUT(n18427));
    defparam add_15136_12.INIT0 = 16'h5aaa;
    defparam add_15136_12.INIT1 = 16'h5aaa;
    defparam add_15136_12.INJECT1_0 = "NO";
    defparam add_15136_12.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i17 (.D(recv_buffer[29]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i18 (.D(recv_buffer[30]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i18.GSR = "DISABLED";
    CCU2D add_15136_10 (.A0(recv_buffer[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18425), .COUT(n18426));
    defparam add_15136_10.INIT0 = 16'h5555;
    defparam add_15136_10.INIT1 = 16'h5aaa;
    defparam add_15136_10.INJECT1_0 = "NO";
    defparam add_15136_10.INJECT1_1 = "NO";
    CCU2D add_15136_8 (.A0(recv_buffer[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18424), .COUT(n18425));
    defparam add_15136_8.INIT0 = 16'h5aaa;
    defparam add_15136_8.INIT1 = 16'h5aaa;
    defparam add_15136_8.INJECT1_0 = "NO";
    defparam add_15136_8.INJECT1_1 = "NO";
    CCU2D add_15136_6 (.A0(recv_buffer[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18423), .COUT(n18424));
    defparam add_15136_6.INIT0 = 16'h5555;
    defparam add_15136_6.INIT1 = 16'h5555;
    defparam add_15136_6.INJECT1_0 = "NO";
    defparam add_15136_6.INJECT1_1 = "NO";
    LUT4 i2763_1_lut (.A(MISO_N_817), .Z(n5199)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(64[1] 216[13])
    defparam i2763_1_lut.init = 16'h5555;
    FD1P3IX speed_set_m1_i0_i1 (.D(recv_buffer[76]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i2 (.D(recv_buffer[77]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i3 (.D(recv_buffer[78]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i4 (.D(recv_buffer[79]), .SP(clkout_c_enable_348), 
            .PD(n14278), .CK(clkout_c), .Q(speed_set_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i5 (.D(recv_buffer[80]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i6 (.D(recv_buffer[81]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i7 (.D(recv_buffer[82]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i8 (.D(recv_buffer[83]), .SP(clkout_c_enable_348), 
            .PD(n14278), .CK(clkout_c), .Q(speed_set_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i9 (.D(recv_buffer[84]), .SP(clkout_c_enable_348), 
            .PD(n14278), .CK(clkout_c), .Q(speed_set_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i9.GSR = "DISABLED";
    CCU2D add_15136_4 (.A0(recv_buffer[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18422), .COUT(n18423));
    defparam add_15136_4.INIT0 = 16'h5aaa;
    defparam add_15136_4.INIT1 = 16'h5555;
    defparam add_15136_4.INJECT1_0 = "NO";
    defparam add_15136_4.INJECT1_1 = "NO";
    FD1P3JX speed_set_m1_i0_i10 (.D(recv_buffer[85]), .SP(clkout_c_enable_348), 
            .PD(n14278), .CK(clkout_c), .Q(speed_set_m1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i11 (.D(recv_buffer[86]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i11.GSR = "DISABLED";
    CCU2D add_15136_2 (.A0(recv_buffer[17]), .B0(recv_buffer[16]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18422));
    defparam add_15136_2.INIT0 = 16'h7000;
    defparam add_15136_2.INIT1 = 16'h5aaa;
    defparam add_15136_2.INJECT1_0 = "NO";
    defparam add_15136_2.INJECT1_1 = "NO";
    FD1P3IX speed_set_m1_i0_i12 (.D(recv_buffer[87]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m1_i0_i13 (.D(recv_buffer[88]), .SP(clkout_c_enable_348), 
            .PD(n14278), .CK(clkout_c), .Q(speed_set_m1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i14 (.D(recv_buffer[89]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i15 (.D(recv_buffer[90]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i16 (.D(recv_buffer[91]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i17 (.D(recv_buffer[92]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i18 (.D(recv_buffer[93]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i19 (.D(recv_buffer[94]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m1_i0_i20 (.D(recv_buffer[95]), .SP(clkout_c_enable_348), 
            .CD(n14278), .CK(clkout_c), .Q(speed_set_m1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m1_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i1 (.D(recv_buffer[55]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i2 (.D(recv_buffer[56]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i3 (.D(recv_buffer[57]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i4 (.D(recv_buffer[58]), .SP(clkout_c_enable_348), 
            .PD(n14258), .CK(clkout_c), .Q(speed_set_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i5 (.D(recv_buffer[59]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i6 (.D(recv_buffer[60]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i7 (.D(recv_buffer[61]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i8 (.D(recv_buffer[62]), .SP(clkout_c_enable_348), 
            .PD(n14258), .CK(clkout_c), .Q(speed_set_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i9 (.D(recv_buffer[63]), .SP(clkout_c_enable_348), 
            .PD(n14258), .CK(clkout_c), .Q(speed_set_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i10 (.D(recv_buffer[64]), .SP(clkout_c_enable_348), 
            .PD(n14258), .CK(clkout_c), .Q(speed_set_m2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i11 (.D(recv_buffer[65]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i12 (.D(recv_buffer[66]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m2_i0_i13 (.D(recv_buffer[67]), .SP(clkout_c_enable_348), 
            .PD(n14258), .CK(clkout_c), .Q(speed_set_m2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i14 (.D(recv_buffer[68]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i15 (.D(recv_buffer[69]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i16 (.D(recv_buffer[70]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i17 (.D(recv_buffer[71]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i18 (.D(recv_buffer[72]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i19 (.D(recv_buffer[73]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m2_i0_i20 (.D(recv_buffer[74]), .SP(clkout_c_enable_348), 
            .CD(n14258), .CK(clkout_c), .Q(speed_set_m2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m2_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i1 (.D(recv_buffer[34]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i1.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i2 (.D(recv_buffer[35]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i3 (.D(recv_buffer[36]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i4 (.D(recv_buffer[37]), .SP(clkout_c_enable_348), 
            .PD(n14238), .CK(clkout_c), .Q(speed_set_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i5 (.D(recv_buffer[38]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i6 (.D(recv_buffer[39]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i7 (.D(recv_buffer[40]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i8 (.D(recv_buffer[41]), .SP(clkout_c_enable_348), 
            .PD(n14238), .CK(clkout_c), .Q(speed_set_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i9 (.D(recv_buffer[42]), .SP(clkout_c_enable_348), 
            .PD(n14238), .CK(clkout_c), .Q(speed_set_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i9.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i10 (.D(recv_buffer[43]), .SP(clkout_c_enable_348), 
            .PD(n14238), .CK(clkout_c), .Q(speed_set_m3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i10.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i11 (.D(recv_buffer[44]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i12 (.D(recv_buffer[45]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m3_i0_i13 (.D(recv_buffer[46]), .SP(clkout_c_enable_348), 
            .PD(n14238), .CK(clkout_c), .Q(speed_set_m3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i13.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i14 (.D(recv_buffer[47]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i14.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i15 (.D(recv_buffer[48]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i15.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i16 (.D(recv_buffer[49]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i16.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i17 (.D(recv_buffer[50]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i17.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i18 (.D(recv_buffer[51]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i18.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i19 (.D(recv_buffer[52]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i20 (.D(recv_buffer[53]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i1 (.D(recv_buffer[13]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i1.GSR = "DISABLED";
    CCU2D add_15139_21 (.A0(recv_buffer[32]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18623), .S1(n3468));
    defparam add_15139_21.INIT0 = 16'h5555;
    defparam add_15139_21.INIT1 = 16'h0000;
    defparam add_15139_21.INJECT1_0 = "NO";
    defparam add_15139_21.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i2 (.D(recv_buffer[14]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i2.GSR = "DISABLED";
    CCU2D add_15139_19 (.A0(recv_buffer[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18622), .COUT(n18623));
    defparam add_15139_19.INIT0 = 16'hf555;
    defparam add_15139_19.INIT1 = 16'hf555;
    defparam add_15139_19.INJECT1_0 = "NO";
    defparam add_15139_19.INJECT1_1 = "NO";
    CCU2D add_15139_17 (.A0(recv_buffer[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18621), .COUT(n18622));
    defparam add_15139_17.INIT0 = 16'hf555;
    defparam add_15139_17.INIT1 = 16'hf555;
    defparam add_15139_17.INJECT1_0 = "NO";
    defparam add_15139_17.INJECT1_1 = "NO";
    CCU2D add_15139_15 (.A0(recv_buffer[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18620), .COUT(n18621));
    defparam add_15139_15.INIT0 = 16'hf555;
    defparam add_15139_15.INIT1 = 16'hf555;
    defparam add_15139_15.INJECT1_0 = "NO";
    defparam add_15139_15.INJECT1_1 = "NO";
    CCU2D add_15139_13 (.A0(recv_buffer[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18619), .COUT(n18620));
    defparam add_15139_13.INIT0 = 16'hf555;
    defparam add_15139_13.INIT1 = 16'h0aaa;
    defparam add_15139_13.INJECT1_0 = "NO";
    defparam add_15139_13.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i3 (.D(recv_buffer[15]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i3.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i4 (.D(recv_buffer[16]), .SP(clkout_c_enable_348), 
            .PD(n14218), .CK(clkout_c), .Q(speed_set_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i4.GSR = "DISABLED";
    CCU2D add_15139_11 (.A0(recv_buffer[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18618), .COUT(n18619));
    defparam add_15139_11.INIT0 = 16'h0aaa;
    defparam add_15139_11.INIT1 = 16'hf555;
    defparam add_15139_11.INJECT1_0 = "NO";
    defparam add_15139_11.INJECT1_1 = "NO";
    CCU2D add_15143_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18479), 
          .S0(n3444));
    defparam add_15143_cout.INIT0 = 16'h0000;
    defparam add_15143_cout.INIT1 = 16'h0000;
    defparam add_15143_cout.INJECT1_0 = "NO";
    defparam add_15143_cout.INJECT1_1 = "NO";
    CCU2D add_15139_9 (.A0(recv_buffer[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18617), .COUT(n18618));
    defparam add_15139_9.INIT0 = 16'h0aaa;
    defparam add_15139_9.INIT1 = 16'h0aaa;
    defparam add_15139_9.INJECT1_0 = "NO";
    defparam add_15139_9.INJECT1_1 = "NO";
    CCU2D add_15139_7 (.A0(recv_buffer[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18616), .COUT(n18617));
    defparam add_15139_7.INIT0 = 16'hf555;
    defparam add_15139_7.INIT1 = 16'hf555;
    defparam add_15139_7.INJECT1_0 = "NO";
    defparam add_15139_7.INJECT1_1 = "NO";
    CCU2D add_15139_5 (.A0(recv_buffer[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18615), .COUT(n18616));
    defparam add_15139_5.INIT0 = 16'h0aaa;
    defparam add_15139_5.INIT1 = 16'hf555;
    defparam add_15139_5.INJECT1_0 = "NO";
    defparam add_15139_5.INJECT1_1 = "NO";
    CCU2D add_15139_3 (.A0(recv_buffer[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18614), .COUT(n18615));
    defparam add_15139_3.INIT0 = 16'hf555;
    defparam add_15139_3.INIT1 = 16'hf555;
    defparam add_15139_3.INJECT1_0 = "NO";
    defparam add_15139_3.INJECT1_1 = "NO";
    CCU2D add_15139_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[12]), .B1(recv_buffer[13]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18614));
    defparam add_15139_1.INIT0 = 16'hF000;
    defparam add_15139_1.INIT1 = 16'ha666;
    defparam add_15139_1.INJECT1_0 = "NO";
    defparam add_15139_1.INJECT1_1 = "NO";
    CCU2D add_15140_21 (.A0(recv_buffer[53]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18603), .S1(n3420));
    defparam add_15140_21.INIT0 = 16'h5555;
    defparam add_15140_21.INIT1 = 16'h0000;
    defparam add_15140_21.INJECT1_0 = "NO";
    defparam add_15140_21.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_388 (.A(CSlatched), .B(CSold), .C(n22211), .Z(clkout_c_enable_348)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i2_3_lut_rep_388.init = 16'h8080;
    LUT4 i11650_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22211), .D(enable_m3_N_834), 
         .Z(n14238)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11650_2_lut_4_lut.init = 16'h0080;
    LUT4 i11690_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22211), .D(enable_m1_N_819), 
         .Z(n14278)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11690_2_lut_4_lut.init = 16'h0080;
    CCU2D add_15140_19 (.A0(recv_buffer[51]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[52]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18602), .COUT(n18603));
    defparam add_15140_19.INIT0 = 16'hf555;
    defparam add_15140_19.INIT1 = 16'hf555;
    defparam add_15140_19.INJECT1_0 = "NO";
    defparam add_15140_19.INJECT1_1 = "NO";
    CCU2D add_15140_17 (.A0(recv_buffer[49]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[50]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18601), .COUT(n18602));
    defparam add_15140_17.INIT0 = 16'hf555;
    defparam add_15140_17.INIT1 = 16'hf555;
    defparam add_15140_17.INJECT1_0 = "NO";
    defparam add_15140_17.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i5 (.D(recv_buffer[17]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i5.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i6 (.D(recv_buffer[18]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i6.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i7 (.D(recv_buffer[19]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i7.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i8 (.D(recv_buffer[20]), .SP(clkout_c_enable_348), 
            .PD(n14218), .CK(clkout_c), .Q(speed_set_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i8.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i9 (.D(recv_buffer[21]), .SP(clkout_c_enable_348), 
            .PD(n14218), .CK(clkout_c), .Q(speed_set_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i9.GSR = "DISABLED";
    CCU2D add_15140_15 (.A0(recv_buffer[47]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[48]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18600), .COUT(n18601));
    defparam add_15140_15.INIT0 = 16'hf555;
    defparam add_15140_15.INIT1 = 16'hf555;
    defparam add_15140_15.INJECT1_0 = "NO";
    defparam add_15140_15.INJECT1_1 = "NO";
    CCU2D add_15140_13 (.A0(recv_buffer[45]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[46]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18599), .COUT(n18600));
    defparam add_15140_13.INIT0 = 16'hf555;
    defparam add_15140_13.INIT1 = 16'h0aaa;
    defparam add_15140_13.INJECT1_0 = "NO";
    defparam add_15140_13.INJECT1_1 = "NO";
    CCU2D add_15140_11 (.A0(recv_buffer[43]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[44]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18598), .COUT(n18599));
    defparam add_15140_11.INIT0 = 16'h0aaa;
    defparam add_15140_11.INIT1 = 16'hf555;
    defparam add_15140_11.INJECT1_0 = "NO";
    defparam add_15140_11.INJECT1_1 = "NO";
    FD1P3JX speed_set_m4_i0_i10 (.D(recv_buffer[22]), .SP(clkout_c_enable_348), 
            .PD(n14218), .CK(clkout_c), .Q(speed_set_m4[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i10.GSR = "DISABLED";
    CCU2D add_15140_9 (.A0(recv_buffer[41]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[42]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18597), .COUT(n18598));
    defparam add_15140_9.INIT0 = 16'h0aaa;
    defparam add_15140_9.INIT1 = 16'h0aaa;
    defparam add_15140_9.INJECT1_0 = "NO";
    defparam add_15140_9.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i11 (.D(recv_buffer[23]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i11.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i12 (.D(recv_buffer[24]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i12.GSR = "DISABLED";
    FD1P3JX speed_set_m4_i0_i13 (.D(recv_buffer[25]), .SP(clkout_c_enable_348), 
            .PD(n14218), .CK(clkout_c), .Q(speed_set_m4[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i13.GSR = "DISABLED";
    CCU2D add_15140_7 (.A0(recv_buffer[39]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[40]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18596), .COUT(n18597));
    defparam add_15140_7.INIT0 = 16'hf555;
    defparam add_15140_7.INIT1 = 16'hf555;
    defparam add_15140_7.INJECT1_0 = "NO";
    defparam add_15140_7.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i14 (.D(recv_buffer[26]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i14.GSR = "DISABLED";
    LUT4 i11630_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22211), .D(enable_m4_N_841), 
         .Z(n14218)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11630_2_lut_4_lut.init = 16'h0080;
    LUT4 i11670_2_lut_4_lut (.A(CSlatched), .B(CSold), .C(n22211), .D(enable_m2_N_827), 
         .Z(n14258)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(139[7:42])
    defparam i11670_2_lut_4_lut.init = 16'h0080;
    CCU2D add_15140_5 (.A0(recv_buffer[37]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[38]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18595), .COUT(n18596));
    defparam add_15140_5.INIT0 = 16'h0aaa;
    defparam add_15140_5.INIT1 = 16'hf555;
    defparam add_15140_5.INJECT1_0 = "NO";
    defparam add_15140_5.INJECT1_1 = "NO";
    CCU2D add_15140_3 (.A0(recv_buffer[35]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[36]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18594), .COUT(n18595));
    defparam add_15140_3.INIT0 = 16'hf555;
    defparam add_15140_3.INIT1 = 16'hf555;
    defparam add_15140_3.INJECT1_0 = "NO";
    defparam add_15140_3.INJECT1_1 = "NO";
    CCU2D add_15140_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[33]), .B1(recv_buffer[34]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18594));
    defparam add_15140_1.INIT0 = 16'hF000;
    defparam add_15140_1.INIT1 = 16'ha666;
    defparam add_15140_1.INJECT1_0 = "NO";
    defparam add_15140_1.INJECT1_1 = "NO";
    FD1P3IX speed_set_m4_i0_i19 (.D(recv_buffer[31]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i19.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i0 (.D(recv_buffer[12]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i0.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i20 (.D(recv_buffer[32]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i20.GSR = "DISABLED";
    FD1P3IX speed_set_m3_i0_i0 (.D(recv_buffer[33]), .SP(clkout_c_enable_348), 
            .CD(n14238), .CK(clkout_c), .Q(speed_set_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m3_i0_i0.GSR = "DISABLED";
    FD1P3IX speed_set_m4_i0_i15 (.D(recv_buffer[27]), .SP(clkout_c_enable_348), 
            .CD(n14218), .CK(clkout_c), .Q(speed_set_m4[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam speed_set_m4_i0_i15.GSR = "DISABLED";
    CCU2D add_15123_21 (.A0(recv_buffer[95]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18570), .S1(n3324));
    defparam add_15123_21.INIT0 = 16'h5555;
    defparam add_15123_21.INIT1 = 16'h0000;
    defparam add_15123_21.INJECT1_0 = "NO";
    defparam add_15123_21.INJECT1_1 = "NO";
    CCU2D add_15123_19 (.A0(recv_buffer[93]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[94]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18569), .COUT(n18570));
    defparam add_15123_19.INIT0 = 16'hf555;
    defparam add_15123_19.INIT1 = 16'hf555;
    defparam add_15123_19.INJECT1_0 = "NO";
    defparam add_15123_19.INJECT1_1 = "NO";
    CCU2D add_15123_17 (.A0(recv_buffer[91]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[92]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18568), .COUT(n18569));
    defparam add_15123_17.INIT0 = 16'hf555;
    defparam add_15123_17.INIT1 = 16'hf555;
    defparam add_15123_17.INJECT1_0 = "NO";
    defparam add_15123_17.INJECT1_1 = "NO";
    CCU2D add_15123_15 (.A0(recv_buffer[89]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[90]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18567), .COUT(n18568));
    defparam add_15123_15.INIT0 = 16'hf555;
    defparam add_15123_15.INIT1 = 16'hf555;
    defparam add_15123_15.INJECT1_0 = "NO";
    defparam add_15123_15.INJECT1_1 = "NO";
    CCU2D add_15123_13 (.A0(recv_buffer[87]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[88]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18566), .COUT(n18567));
    defparam add_15123_13.INIT0 = 16'hf555;
    defparam add_15123_13.INIT1 = 16'h0aaa;
    defparam add_15123_13.INJECT1_0 = "NO";
    defparam add_15123_13.INJECT1_1 = "NO";
    CCU2D add_15123_11 (.A0(recv_buffer[85]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[86]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18565), .COUT(n18566));
    defparam add_15123_11.INIT0 = 16'h0aaa;
    defparam add_15123_11.INIT1 = 16'hf555;
    defparam add_15123_11.INJECT1_0 = "NO";
    defparam add_15123_11.INJECT1_1 = "NO";
    CCU2D add_15123_9 (.A0(recv_buffer[83]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[84]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18564), .COUT(n18565));
    defparam add_15123_9.INIT0 = 16'h0aaa;
    defparam add_15123_9.INIT1 = 16'h0aaa;
    defparam add_15123_9.INJECT1_0 = "NO";
    defparam add_15123_9.INJECT1_1 = "NO";
    CCU2D add_15123_7 (.A0(recv_buffer[81]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[82]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18563), .COUT(n18564));
    defparam add_15123_7.INIT0 = 16'hf555;
    defparam add_15123_7.INIT1 = 16'hf555;
    defparam add_15123_7.INJECT1_0 = "NO";
    defparam add_15123_7.INJECT1_1 = "NO";
    CCU2D add_15123_5 (.A0(recv_buffer[79]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[80]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18562), .COUT(n18563));
    defparam add_15123_5.INIT0 = 16'h0aaa;
    defparam add_15123_5.INIT1 = 16'hf555;
    defparam add_15123_5.INJECT1_0 = "NO";
    defparam add_15123_5.INJECT1_1 = "NO";
    CCU2D add_15123_3 (.A0(recv_buffer[77]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[78]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18561), .COUT(n18562));
    defparam add_15123_3.INIT0 = 16'hf555;
    defparam add_15123_3.INIT1 = 16'hf555;
    defparam add_15123_3.INJECT1_0 = "NO";
    defparam add_15123_3.INJECT1_1 = "NO";
    CCU2D add_15123_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(recv_buffer[75]), .B1(recv_buffer[76]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18561));
    defparam add_15123_1.INIT0 = 16'hF000;
    defparam add_15123_1.INIT1 = 16'ha666;
    defparam add_15123_1.INJECT1_0 = "NO";
    defparam add_15123_1.INJECT1_1 = "NO";
    CCU2D add_15141_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18560), 
          .S0(n3396));
    defparam add_15141_cout.INIT0 = 16'h0000;
    defparam add_15141_cout.INIT1 = 16'h0000;
    defparam add_15141_cout.INJECT1_0 = "NO";
    defparam add_15141_cout.INJECT1_1 = "NO";
    CCU2D add_15141_16 (.A0(recv_buffer[73]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[74]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18559), .COUT(n18560));
    defparam add_15141_16.INIT0 = 16'h5aaa;
    defparam add_15141_16.INIT1 = 16'h0aaa;
    defparam add_15141_16.INJECT1_0 = "NO";
    defparam add_15141_16.INJECT1_1 = "NO";
    CCU2D add_15141_14 (.A0(recv_buffer[71]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[72]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18558), .COUT(n18559));
    defparam add_15141_14.INIT0 = 16'h5aaa;
    defparam add_15141_14.INIT1 = 16'h5aaa;
    defparam add_15141_14.INJECT1_0 = "NO";
    defparam add_15141_14.INJECT1_1 = "NO";
    CCU2D add_15141_12 (.A0(recv_buffer[69]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[70]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18557), .COUT(n18558));
    defparam add_15141_12.INIT0 = 16'h5aaa;
    defparam add_15141_12.INIT1 = 16'h5aaa;
    defparam add_15141_12.INJECT1_0 = "NO";
    defparam add_15141_12.INJECT1_1 = "NO";
    CCU2D add_15141_10 (.A0(recv_buffer[67]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[68]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18556), .COUT(n18557));
    defparam add_15141_10.INIT0 = 16'h5555;
    defparam add_15141_10.INIT1 = 16'h5aaa;
    defparam add_15141_10.INJECT1_0 = "NO";
    defparam add_15141_10.INJECT1_1 = "NO";
    CCU2D add_15141_8 (.A0(recv_buffer[65]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[66]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18555), .COUT(n18556));
    defparam add_15141_8.INIT0 = 16'h5aaa;
    defparam add_15141_8.INIT1 = 16'h5aaa;
    defparam add_15141_8.INJECT1_0 = "NO";
    defparam add_15141_8.INJECT1_1 = "NO";
    CCU2D add_15141_6 (.A0(recv_buffer[63]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[64]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18554), .COUT(n18555));
    defparam add_15141_6.INIT0 = 16'h5555;
    defparam add_15141_6.INIT1 = 16'h5555;
    defparam add_15141_6.INJECT1_0 = "NO";
    defparam add_15141_6.INJECT1_1 = "NO";
    CCU2D add_15141_4 (.A0(recv_buffer[61]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[62]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18553), .COUT(n18554));
    defparam add_15141_4.INIT0 = 16'h5aaa;
    defparam add_15141_4.INIT1 = 16'h5555;
    defparam add_15141_4.INJECT1_0 = "NO";
    defparam add_15141_4.INJECT1_1 = "NO";
    CCU2D add_15141_2 (.A0(recv_buffer[59]), .B0(recv_buffer[58]), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[60]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18553));
    defparam add_15141_2.INIT0 = 16'h7000;
    defparam add_15141_2.INIT1 = 16'h5aaa;
    defparam add_15141_2.INJECT1_0 = "NO";
    defparam add_15141_2.INJECT1_1 = "NO";
    CCU2D add_15143_16 (.A0(recv_buffer[52]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[53]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18478), .COUT(n18479));
    defparam add_15143_16.INIT0 = 16'h5aaa;
    defparam add_15143_16.INIT1 = 16'h0aaa;
    defparam add_15143_16.INJECT1_0 = "NO";
    defparam add_15143_16.INJECT1_1 = "NO";
    CCU2D add_15143_14 (.A0(recv_buffer[50]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[51]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18477), .COUT(n18478));
    defparam add_15143_14.INIT0 = 16'h5aaa;
    defparam add_15143_14.INIT1 = 16'h5aaa;
    defparam add_15143_14.INJECT1_0 = "NO";
    defparam add_15143_14.INJECT1_1 = "NO";
    CCU2D add_15143_12 (.A0(recv_buffer[48]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(recv_buffer[49]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18476), .COUT(n18477));
    defparam add_15143_12.INIT0 = 16'h5aaa;
    defparam add_15143_12.INIT1 = 16'h5aaa;
    defparam add_15143_12.INJECT1_0 = "NO";
    defparam add_15143_12.INJECT1_1 = "NO";
    FD1P3AX CSold_116_rep_402 (.D(n22207), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(n22208));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSold_116_rep_402.GSR = "DISABLED";
    FD1P3AX CSlatched_118_rep_401 (.D(CS_c), .SP(clkout_c_enable_362), .CK(clkout_c), 
            .Q(n22207));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/spi loopbacktest v2.vhd(89[2] 213[9])
    defparam CSlatched_118_rep_401.GSR = "DISABLED";
    PFUMX MISO_I_0 (.BLUT(n5197), .ALUT(MISOb_N_857), .C0(n22211), .Z(MISO_N_862)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=313, LSE_RLINE=313 */ ;
    
endmodule
//
// Verilog Description of module AVG_SPEED_U9
//

module AVG_SPEED_U9 (\speed_avg_m3[0] , clk_1mhz, \speed_m3[0] , \speed_avg_m3[1] , 
            \speed_m3[1] , \speed_avg_m3[2] , \speed_m3[2] , \speed_avg_m3[3] , 
            \speed_m3[3] , \speed_avg_m3[4] , \speed_m3[4] , \speed_avg_m3[5] , 
            \speed_m3[5] , \speed_avg_m3[6] , \speed_m3[6] , \speed_avg_m3[7] , 
            \speed_m3[7] , \speed_avg_m3[8] , \speed_m3[8] , \speed_avg_m3[9] , 
            \speed_m3[9] , \speed_avg_m3[10] , \speed_m3[10] , \speed_avg_m3[11] , 
            \speed_m3[11] , \speed_avg_m3[12] , \speed_m3[12] , \speed_avg_m3[13] , 
            \speed_m3[13] , \speed_avg_m3[14] , \speed_m3[14] , \speed_avg_m3[15] , 
            \speed_m3[15] , \speed_avg_m3[16] , \speed_m3[16] , \speed_avg_m3[17] , 
            \speed_m3[17] , \speed_avg_m3[18] , \speed_m3[18] , \speed_avg_m3[19] , 
            \speed_m3[19] , GND_net);
    output \speed_avg_m3[0] ;
    input clk_1mhz;
    input \speed_m3[0] ;
    output \speed_avg_m3[1] ;
    input \speed_m3[1] ;
    output \speed_avg_m3[2] ;
    input \speed_m3[2] ;
    output \speed_avg_m3[3] ;
    input \speed_m3[3] ;
    output \speed_avg_m3[4] ;
    input \speed_m3[4] ;
    output \speed_avg_m3[5] ;
    input \speed_m3[5] ;
    output \speed_avg_m3[6] ;
    input \speed_m3[6] ;
    output \speed_avg_m3[7] ;
    input \speed_m3[7] ;
    output \speed_avg_m3[8] ;
    input \speed_m3[8] ;
    output \speed_avg_m3[9] ;
    input \speed_m3[9] ;
    output \speed_avg_m3[10] ;
    input \speed_m3[10] ;
    output \speed_avg_m3[11] ;
    input \speed_m3[11] ;
    output \speed_avg_m3[12] ;
    input \speed_m3[12] ;
    output \speed_avg_m3[13] ;
    input \speed_m3[13] ;
    output \speed_avg_m3[14] ;
    input \speed_m3[14] ;
    output \speed_avg_m3[15] ;
    input \speed_m3[15] ;
    output \speed_avg_m3[16] ;
    input \speed_m3[16] ;
    output \speed_avg_m3[17] ;
    input \speed_m3[17] ;
    output \speed_avg_m3[18] ;
    input \speed_m3[18] ;
    output \speed_avg_m3[19] ;
    input \speed_m3[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_145;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n19871, n6, n18377, n18376, n18375;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m3[0] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2136__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_145), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136__i0.GSR = "DISABLED";
    LUT4 i17245_4_lut (.A(clk_cnt[4]), .B(n19871), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_145)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17245_4_lut.init = 16'h0004;
    LUT4 i16419_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n19871)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16419_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i1_2_lut.init = 16'heeee;
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m3[1] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m3[2] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m3[3] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m3[4] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m3[5] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m3[6] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m3[7] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m3[8] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m3[9] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m3[10] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m3[11] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m3[12] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m3[13] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m3[14] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m3[15] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m3[16] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m3[17] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m3[18] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m3[19] ), .SP(clk_1mhz_enable_145), 
            .CK(clk_1mhz), .Q(\speed_avg_m3[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=367, LSE_RLINE=367 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    CCU2D clk_cnt_2136_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18377), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2136_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2136_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2136_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2136_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18376), .COUT(n18377), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2136_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2136_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2136_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2136_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18375), .COUT(n18376), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2136_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2136_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2136_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2136_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18375), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2136_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2136_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2136_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2136__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_145), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2136__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_145), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2136__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_145), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2136__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_145), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2136__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_145), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2136__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_145), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2136__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module AVG_SPEED_U10
//

module AVG_SPEED_U10 (\speed_avg_m2[0] , clk_1mhz, \speed_m2[0] , \speed_avg_m2[1] , 
            \speed_m2[1] , \speed_avg_m2[2] , \speed_m2[2] , \speed_avg_m2[3] , 
            \speed_m2[3] , \speed_avg_m2[4] , \speed_m2[4] , \speed_avg_m2[5] , 
            \speed_m2[5] , \speed_avg_m2[6] , \speed_m2[6] , \speed_avg_m2[7] , 
            \speed_m2[7] , \speed_avg_m2[8] , \speed_m2[8] , \speed_avg_m2[9] , 
            \speed_m2[9] , \speed_avg_m2[10] , \speed_m2[10] , \speed_avg_m2[11] , 
            \speed_m2[11] , \speed_avg_m2[12] , \speed_m2[12] , \speed_avg_m2[13] , 
            \speed_m2[13] , \speed_avg_m2[14] , \speed_m2[14] , \speed_avg_m2[15] , 
            \speed_m2[15] , \speed_avg_m2[16] , \speed_m2[16] , \speed_avg_m2[17] , 
            \speed_m2[17] , \speed_avg_m2[18] , \speed_m2[18] , \speed_avg_m2[19] , 
            \speed_m2[19] , GND_net);
    output \speed_avg_m2[0] ;
    input clk_1mhz;
    input \speed_m2[0] ;
    output \speed_avg_m2[1] ;
    input \speed_m2[1] ;
    output \speed_avg_m2[2] ;
    input \speed_m2[2] ;
    output \speed_avg_m2[3] ;
    input \speed_m2[3] ;
    output \speed_avg_m2[4] ;
    input \speed_m2[4] ;
    output \speed_avg_m2[5] ;
    input \speed_m2[5] ;
    output \speed_avg_m2[6] ;
    input \speed_m2[6] ;
    output \speed_avg_m2[7] ;
    input \speed_m2[7] ;
    output \speed_avg_m2[8] ;
    input \speed_m2[8] ;
    output \speed_avg_m2[9] ;
    input \speed_m2[9] ;
    output \speed_avg_m2[10] ;
    input \speed_m2[10] ;
    output \speed_avg_m2[11] ;
    input \speed_m2[11] ;
    output \speed_avg_m2[12] ;
    input \speed_m2[12] ;
    output \speed_avg_m2[13] ;
    input \speed_m2[13] ;
    output \speed_avg_m2[14] ;
    input \speed_m2[14] ;
    output \speed_avg_m2[15] ;
    input \speed_m2[15] ;
    output \speed_avg_m2[16] ;
    input \speed_m2[16] ;
    output \speed_avg_m2[17] ;
    input \speed_m2[17] ;
    output \speed_avg_m2[18] ;
    input \speed_m2[18] ;
    output \speed_avg_m2[19] ;
    input \speed_m2[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_126;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n19849, n6, n18381, n18380, n18379;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m2[0] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2134__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_126), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134__i0.GSR = "DISABLED";
    LUT4 i17251_4_lut (.A(clk_cnt[0]), .B(n19849), .C(clk_cnt[3]), .D(n6), 
         .Z(clk_1mhz_enable_126)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17251_4_lut.init = 16'h0004;
    LUT4 i16397_3_lut (.A(clk_cnt[2]), .B(clk_cnt[6]), .C(clk_cnt[5]), 
         .Z(n19849)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16397_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(clk_cnt[1]), .B(clk_cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m2[1] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m2[2] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m2[3] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m2[4] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m2[5] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m2[6] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m2[7] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m2[8] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m2[9] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m2[10] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m2[11] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m2[12] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m2[13] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m2[14] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m2[15] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m2[16] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m2[17] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m2[18] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m2[19] ), .SP(clk_1mhz_enable_126), 
            .CK(clk_1mhz), .Q(\speed_avg_m2[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=364, LSE_RLINE=364 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    CCU2D clk_cnt_2134_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18381), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2134_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2134_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2134_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2134_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18380), .COUT(n18381), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2134_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2134_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2134_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2134_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18379), .COUT(n18380), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2134_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2134_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2134_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2134_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18379), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2134_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2134_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2134_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2134__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_126), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2134__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_126), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2134__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_126), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2134__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_126), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2134__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_126), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2134__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_126), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2134__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module AVG_SPEED_U11
//

module AVG_SPEED_U11 (\speed_avg_m1[0] , clk_1mhz, \speed_m1[0] , \speed_avg_m1[1] , 
            \speed_m1[1] , \speed_avg_m1[2] , \speed_m1[2] , \speed_avg_m1[3] , 
            \speed_m1[3] , \speed_avg_m1[4] , \speed_m1[4] , \speed_avg_m1[5] , 
            \speed_m1[5] , \speed_avg_m1[6] , \speed_m1[6] , \speed_avg_m1[7] , 
            \speed_m1[7] , \speed_avg_m1[8] , \speed_m1[8] , \speed_avg_m1[9] , 
            \speed_m1[9] , \speed_avg_m1[10] , \speed_m1[10] , \speed_avg_m1[11] , 
            \speed_m1[11] , \speed_avg_m1[12] , \speed_m1[12] , \speed_avg_m1[13] , 
            \speed_m1[13] , \speed_avg_m1[14] , \speed_m1[14] , \speed_avg_m1[15] , 
            \speed_m1[15] , \speed_avg_m1[16] , \speed_m1[16] , \speed_avg_m1[17] , 
            \speed_m1[17] , \speed_avg_m1[18] , \speed_m1[18] , \speed_avg_m1[19] , 
            \speed_m1[19] , GND_net);
    output \speed_avg_m1[0] ;
    input clk_1mhz;
    input \speed_m1[0] ;
    output \speed_avg_m1[1] ;
    input \speed_m1[1] ;
    output \speed_avg_m1[2] ;
    input \speed_m1[2] ;
    output \speed_avg_m1[3] ;
    input \speed_m1[3] ;
    output \speed_avg_m1[4] ;
    input \speed_m1[4] ;
    output \speed_avg_m1[5] ;
    input \speed_m1[5] ;
    output \speed_avg_m1[6] ;
    input \speed_m1[6] ;
    output \speed_avg_m1[7] ;
    input \speed_m1[7] ;
    output \speed_avg_m1[8] ;
    input \speed_m1[8] ;
    output \speed_avg_m1[9] ;
    input \speed_m1[9] ;
    output \speed_avg_m1[10] ;
    input \speed_m1[10] ;
    output \speed_avg_m1[11] ;
    input \speed_m1[11] ;
    output \speed_avg_m1[12] ;
    input \speed_m1[12] ;
    output \speed_avg_m1[13] ;
    input \speed_m1[13] ;
    output \speed_avg_m1[14] ;
    input \speed_m1[14] ;
    output \speed_avg_m1[15] ;
    input \speed_m1[15] ;
    output \speed_avg_m1[16] ;
    input \speed_m1[16] ;
    output \speed_avg_m1[17] ;
    input \speed_m1[17] ;
    output \speed_avg_m1[18] ;
    input \speed_m1[18] ;
    output \speed_avg_m1[19] ;
    input \speed_m1[19] ;
    input GND_net;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    
    wire clk_1mhz_enable_107;
    wire [6:0]clk_cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(31[9:16])
    wire [6:0]n33;
    
    wire n12, n18385, n18384, n18383;
    
    FD1P3AX speed_avg_i0_i0 (.D(\speed_m1[0] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i0.GSR = "DISABLED";
    FD1S3IX clk_cnt_2132__i0 (.D(n33[0]), .CK(clk_1mhz), .CD(clk_1mhz_enable_107), 
            .Q(clk_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132__i0.GSR = "DISABLED";
    LUT4 i17248_4_lut (.A(clk_cnt[2]), .B(n12), .C(clk_cnt[1]), .D(clk_cnt[6]), 
         .Z(clk_1mhz_enable_107)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(49[5:18])
    defparam i17248_4_lut.init = 16'h0200;
    LUT4 i5_4_lut (.A(clk_cnt[4]), .B(clk_cnt[3]), .C(clk_cnt[0]), .D(clk_cnt[5]), 
         .Z(n12)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i5_4_lut.init = 16'hfeff;
    FD1P3AX speed_avg_i0_i1 (.D(\speed_m1[1] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i1.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i2 (.D(\speed_m1[2] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i2.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i3 (.D(\speed_m1[3] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i3.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i4 (.D(\speed_m1[4] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i4.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i5 (.D(\speed_m1[5] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i5.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i6 (.D(\speed_m1[6] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i6.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i7 (.D(\speed_m1[7] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i7.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i8 (.D(\speed_m1[8] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i8.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i9 (.D(\speed_m1[9] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i9.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i10 (.D(\speed_m1[10] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i10.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i11 (.D(\speed_m1[11] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i11.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i12 (.D(\speed_m1[12] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i12.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i13 (.D(\speed_m1[13] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i13.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i14 (.D(\speed_m1[14] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i14.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i15 (.D(\speed_m1[15] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i15.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i16 (.D(\speed_m1[16] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i16.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i17 (.D(\speed_m1[17] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i17.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i18 (.D(\speed_m1[18] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i18.GSR = "DISABLED";
    FD1P3AX speed_avg_i0_i19 (.D(\speed_m1[19] ), .SP(clk_1mhz_enable_107), 
            .CK(clk_1mhz), .Q(\speed_avg_m1[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=17, LSE_RCOL=26, LSE_LLINE=361, LSE_RLINE=361 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(46[1] 66[8])
    defparam speed_avg_i0_i19.GSR = "DISABLED";
    CCU2D clk_cnt_2132_add_4_7 (.A0(clk_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18385), .S0(n33[5]), .S1(n33[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132_add_4_7.INIT0 = 16'hfaaa;
    defparam clk_cnt_2132_add_4_7.INIT1 = 16'hfaaa;
    defparam clk_cnt_2132_add_4_7.INJECT1_0 = "NO";
    defparam clk_cnt_2132_add_4_7.INJECT1_1 = "NO";
    CCU2D clk_cnt_2132_add_4_5 (.A0(clk_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18384), .COUT(n18385), .S0(n33[3]), .S1(n33[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132_add_4_5.INIT0 = 16'hfaaa;
    defparam clk_cnt_2132_add_4_5.INIT1 = 16'hfaaa;
    defparam clk_cnt_2132_add_4_5.INJECT1_0 = "NO";
    defparam clk_cnt_2132_add_4_5.INJECT1_1 = "NO";
    CCU2D clk_cnt_2132_add_4_3 (.A0(clk_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18383), .COUT(n18384), .S0(n33[1]), .S1(n33[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132_add_4_3.INIT0 = 16'hfaaa;
    defparam clk_cnt_2132_add_4_3.INIT1 = 16'hfaaa;
    defparam clk_cnt_2132_add_4_3.INJECT1_0 = "NO";
    defparam clk_cnt_2132_add_4_3.INJECT1_1 = "NO";
    CCU2D clk_cnt_2132_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(clk_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18383), .S1(n33[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132_add_4_1.INIT0 = 16'hF000;
    defparam clk_cnt_2132_add_4_1.INIT1 = 16'h0555;
    defparam clk_cnt_2132_add_4_1.INJECT1_0 = "NO";
    defparam clk_cnt_2132_add_4_1.INJECT1_1 = "NO";
    FD1S3IX clk_cnt_2132__i1 (.D(n33[1]), .CK(clk_1mhz), .CD(clk_1mhz_enable_107), 
            .Q(clk_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132__i1.GSR = "DISABLED";
    FD1S3IX clk_cnt_2132__i2 (.D(n33[2]), .CK(clk_1mhz), .CD(clk_1mhz_enable_107), 
            .Q(clk_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132__i2.GSR = "DISABLED";
    FD1S3IX clk_cnt_2132__i3 (.D(n33[3]), .CK(clk_1mhz), .CD(clk_1mhz_enable_107), 
            .Q(clk_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132__i3.GSR = "DISABLED";
    FD1S3IX clk_cnt_2132__i4 (.D(n33[4]), .CK(clk_1mhz), .CD(clk_1mhz_enable_107), 
            .Q(clk_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132__i4.GSR = "DISABLED";
    FD1S3IX clk_cnt_2132__i5 (.D(n33[5]), .CK(clk_1mhz), .CD(clk_1mhz_enable_107), 
            .Q(clk_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132__i5.GSR = "DISABLED";
    FD1S3IX clk_cnt_2132__i6 (.D(n33[6]), .CK(clk_1mhz), .CD(clk_1mhz_enable_107), 
            .Q(clk_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/speed_avg.vhd(62[14:21])
    defparam clk_cnt_2132__i6.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U1
//

module PWMGENERATOR_U1 (PWM_m2, pwm_clk, LED2_c, clkout_c_enable_362, 
            PWMdut_m2, GND_net);
    output PWM_m2;
    input pwm_clk;
    output LED2_c;
    input clkout_c_enable_362;
    input [9:0]PWMdut_m2;
    input GND_net;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire PWM_N_2176, free_N_2188, n3866, n7;
    wire [9:0]n1;
    
    wire n7_adj_2390, n8, n11549, n14, n10_adj_2391, n17;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    
    wire n16, n14215, n18401;
    wire [9:0]n45;
    
    wire n18400, n18399, n18398, n18397, n21436, n18358, n18357, 
        n18356, n18355, n18354;
    
    FD1S3AX PWM_22 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m2)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=338, LSE_RLINE=338 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam PWM_22.GSR = "ENABLED";
    FD1P3AX free_21 (.D(free_N_2188), .SP(clkout_c_enable_362), .CK(pwm_clk), 
            .Q(LED2_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam free_21.GSR = "DISABLED";
    LUT4 i1806_1_lut (.A(n3866), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1806_1_lut.init = 16'h5555;
    LUT4 i13286_2_lut (.A(PWMdut_m2[8]), .B(n7), .Z(n1[8])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13286_2_lut.init = 16'heeee;
    LUT4 i5_4_lut (.A(PWMdut_m2[9]), .B(n7_adj_2390), .C(PWMdut_m2[7]), 
         .D(n8), .Z(n7)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(PWMdut_m2[6]), .B(n11549), .C(PWMdut_m2[4]), .D(PWMdut_m2[3]), 
         .Z(n7_adj_2390)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut.init = 16'ha8a0;
    LUT4 i2_2_lut (.A(PWMdut_m2[5]), .B(PWMdut_m2[8]), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i13284_2_lut (.A(PWMdut_m2[6]), .B(n7), .Z(n1[6])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13284_2_lut.init = 16'heeee;
    LUT4 i13282_2_lut (.A(PWMdut_m2[3]), .B(n7), .Z(n1[3])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13282_2_lut.init = 16'heeee;
    LUT4 i6_4_lut (.A(PWMdut_m2[9]), .B(PWMdut_m2[3]), .C(PWMdut_m2[4]), 
         .D(n11549), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_adj_150 (.A(PWMdut_m2[6]), .B(PWMdut_m2[7]), .Z(n10_adj_2391)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut_adj_150.init = 16'heeee;
    LUT4 i2_3_lut (.A(PWMdut_m2[2]), .B(PWMdut_m2[1]), .C(PWMdut_m2[0]), 
         .Z(n11549)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i17195_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n14215)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(77[6:16])
    defparam i17195_4_lut.init = 16'h0400;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i6_4_lut_adj_151 (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), 
         .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut_adj_151.init = 16'hffef;
    CCU2D cnt_2128_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18401), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2128_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2128_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2128_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2128_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18400), 
          .COUT(n18401), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2128_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2128_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2128_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2128_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18399), 
          .COUT(n18400), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2128_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2128_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2128_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2128_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18398), 
          .COUT(n18399), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2128_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2128_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2128_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2128_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18397), 
          .COUT(n18398), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2128_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2128_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2128_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2128_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18397), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2128_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2128_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2128_add_4_1.INJECT1_1 = "NO";
    LUT4 i7_4_lut_rep_335 (.A(PWMdut_m2[5]), .B(n14), .C(n10_adj_2391), 
         .D(PWMdut_m2[8]), .Z(n21436)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i7_4_lut_rep_335.init = 16'hfffe;
    LUT4 DutyCycle_9__I_0_i20_1_lut_4_lut (.A(PWMdut_m2[5]), .B(n14), .C(n10_adj_2391), 
         .D(PWMdut_m2[8]), .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam DutyCycle_9__I_0_i20_1_lut_4_lut.init = 16'h0001;
    CCU2D sub_1804_add_2_11 (.A0(PWMdut_m2[9]), .B0(n21436), .C0(cnt[9]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18358), .S1(n3866));
    defparam sub_1804_add_2_11.INIT0 = 16'h8787;
    defparam sub_1804_add_2_11.INIT1 = 16'h0000;
    defparam sub_1804_add_2_11.INJECT1_0 = "NO";
    defparam sub_1804_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_9 (.A0(PWMdut_m2[7]), .B0(n21436), .C0(cnt[7]), 
          .D0(GND_net), .A1(n1[8]), .B1(n21436), .C1(cnt[8]), .D1(GND_net), 
          .CIN(n18357), .COUT(n18358));
    defparam sub_1804_add_2_9.INIT0 = 16'h8787;
    defparam sub_1804_add_2_9.INIT1 = 16'h8787;
    defparam sub_1804_add_2_9.INJECT1_0 = "NO";
    defparam sub_1804_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_7 (.A0(PWMdut_m2[5]), .B0(n21436), .C0(cnt[5]), 
          .D0(GND_net), .A1(n1[6]), .B1(n21436), .C1(cnt[6]), .D1(GND_net), 
          .CIN(n18356), .COUT(n18357));
    defparam sub_1804_add_2_7.INIT0 = 16'h8787;
    defparam sub_1804_add_2_7.INIT1 = 16'h8787;
    defparam sub_1804_add_2_7.INJECT1_0 = "NO";
    defparam sub_1804_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_5 (.A0(n1[3]), .B0(n21436), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(n21436), .C1(n7), .D1(PWMdut_m2[4]), .CIN(n18355), 
          .COUT(n18356));
    defparam sub_1804_add_2_5.INIT0 = 16'h8787;
    defparam sub_1804_add_2_5.INIT1 = 16'h5955;
    defparam sub_1804_add_2_5.INJECT1_0 = "NO";
    defparam sub_1804_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_3 (.A0(cnt[1]), .B0(n21436), .C0(n7), .D0(PWMdut_m2[1]), 
          .A1(cnt[2]), .B1(n21436), .C1(n7), .D1(PWMdut_m2[2]), .CIN(n18354), 
          .COUT(n18355));
    defparam sub_1804_add_2_3.INIT0 = 16'h5955;
    defparam sub_1804_add_2_3.INIT1 = 16'h5955;
    defparam sub_1804_add_2_3.INJECT1_0 = "NO";
    defparam sub_1804_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1804_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(n21436), .C1(n7), .D1(PWMdut_m2[0]), 
          .COUT(n18354));
    defparam sub_1804_add_2_1.INIT0 = 16'h0000;
    defparam sub_1804_add_2_1.INIT1 = 16'h5955;
    defparam sub_1804_add_2_1.INJECT1_0 = "NO";
    defparam sub_1804_add_2_1.INJECT1_1 = "NO";
    FD1S3IX cnt_2128__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14215), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i0.GSR = "ENABLED";
    FD1S3IX cnt_2128__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14215), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i1.GSR = "ENABLED";
    FD1S3IX cnt_2128__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14215), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i2.GSR = "ENABLED";
    FD1S3IX cnt_2128__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14215), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i3.GSR = "ENABLED";
    FD1S3IX cnt_2128__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14215), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i4.GSR = "ENABLED";
    FD1S3IX cnt_2128__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14215), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i5.GSR = "ENABLED";
    FD1S3IX cnt_2128__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14215), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i6.GSR = "ENABLED";
    FD1S3IX cnt_2128__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14215), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i7.GSR = "ENABLED";
    FD1S3IX cnt_2128__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14215), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i8.GSR = "ENABLED";
    FD1S3IX cnt_2128__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14215), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2128__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U0
//

module PWMGENERATOR_U0 (PWMdut_m3, GND_net, PWM_m3, pwm_clk, LED3_c, 
            clkout_c_enable_362);
    input [9:0]PWMdut_m3;
    input GND_net;
    output PWM_m3;
    input pwm_clk;
    output LED3_c;
    input clkout_c_enable_362;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire n18343, n21434;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    
    wire n3879, n18342;
    wire [9:0]n1;
    
    wire n18341, n18340, n7, n18339, PWM_N_2176, free_N_2188, n7_adj_2388, 
        n8, n11551, n19915, n6, n14214, n19899, n14, n10_adj_2389, 
        n18396;
    wire [9:0]n45;
    
    wire n18395, n18394, n18393, n18392;
    
    CCU2D sub_1806_add_2_11 (.A0(PWMdut_m3[9]), .B0(n21434), .C0(cnt[9]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18343), .S1(n3879));
    defparam sub_1806_add_2_11.INIT0 = 16'h8787;
    defparam sub_1806_add_2_11.INIT1 = 16'h0000;
    defparam sub_1806_add_2_11.INJECT1_0 = "NO";
    defparam sub_1806_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_9 (.A0(PWMdut_m3[7]), .B0(n21434), .C0(cnt[7]), 
          .D0(GND_net), .A1(n1[8]), .B1(n21434), .C1(cnt[8]), .D1(GND_net), 
          .CIN(n18342), .COUT(n18343));
    defparam sub_1806_add_2_9.INIT0 = 16'h8787;
    defparam sub_1806_add_2_9.INIT1 = 16'h8787;
    defparam sub_1806_add_2_9.INJECT1_0 = "NO";
    defparam sub_1806_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_7 (.A0(PWMdut_m3[5]), .B0(n21434), .C0(cnt[5]), 
          .D0(GND_net), .A1(n1[6]), .B1(n21434), .C1(cnt[6]), .D1(GND_net), 
          .CIN(n18341), .COUT(n18342));
    defparam sub_1806_add_2_7.INIT0 = 16'h8787;
    defparam sub_1806_add_2_7.INIT1 = 16'h8787;
    defparam sub_1806_add_2_7.INJECT1_0 = "NO";
    defparam sub_1806_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_5 (.A0(n1[3]), .B0(n21434), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(n21434), .C1(n7), .D1(PWMdut_m3[4]), .CIN(n18340), 
          .COUT(n18341));
    defparam sub_1806_add_2_5.INIT0 = 16'h8787;
    defparam sub_1806_add_2_5.INIT1 = 16'h5955;
    defparam sub_1806_add_2_5.INJECT1_0 = "NO";
    defparam sub_1806_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_3 (.A0(cnt[1]), .B0(n21434), .C0(n7), .D0(PWMdut_m3[1]), 
          .A1(cnt[2]), .B1(n21434), .C1(n7), .D1(PWMdut_m3[2]), .CIN(n18339), 
          .COUT(n18340));
    defparam sub_1806_add_2_3.INIT0 = 16'h5955;
    defparam sub_1806_add_2_3.INIT1 = 16'h5955;
    defparam sub_1806_add_2_3.INJECT1_0 = "NO";
    defparam sub_1806_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1806_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(n21434), .C1(n7), .D1(PWMdut_m3[0]), 
          .COUT(n18339));
    defparam sub_1806_add_2_1.INIT0 = 16'h0000;
    defparam sub_1806_add_2_1.INIT1 = 16'h5955;
    defparam sub_1806_add_2_1.INJECT1_0 = "NO";
    defparam sub_1806_add_2_1.INJECT1_1 = "NO";
    FD1S3AX PWM_22 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m3)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=348, LSE_RLINE=348 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam PWM_22.GSR = "ENABLED";
    FD1P3AX free_21 (.D(free_N_2188), .SP(clkout_c_enable_362), .CK(pwm_clk), 
            .Q(LED3_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam free_21.GSR = "DISABLED";
    LUT4 i13303_2_lut (.A(PWMdut_m3[8]), .B(n7), .Z(n1[8])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13303_2_lut.init = 16'heeee;
    LUT4 i5_4_lut (.A(PWMdut_m3[9]), .B(n7_adj_2388), .C(PWMdut_m3[7]), 
         .D(n8), .Z(n7)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(PWMdut_m3[6]), .B(n11551), .C(PWMdut_m3[4]), .D(PWMdut_m3[3]), 
         .Z(n7_adj_2388)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut.init = 16'ha8a0;
    LUT4 i2_2_lut (.A(PWMdut_m3[5]), .B(PWMdut_m3[8]), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i13301_2_lut (.A(PWMdut_m3[6]), .B(n7), .Z(n1[6])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13301_2_lut.init = 16'heeee;
    LUT4 i13299_2_lut (.A(PWMdut_m3[3]), .B(n7), .Z(n1[3])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13299_2_lut.init = 16'heeee;
    LUT4 i1808_1_lut (.A(n3879), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1808_1_lut.init = 16'h5555;
    LUT4 i17192_4_lut (.A(cnt[0]), .B(n19915), .C(cnt[2]), .D(n6), .Z(n14214)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(77[6:16])
    defparam i17192_4_lut.init = 16'h0004;
    LUT4 i16463_3_lut (.A(cnt[7]), .B(n19899), .C(cnt[3]), .Z(n19915)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16463_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[1]), .B(cnt[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i16447_4_lut (.A(cnt[8]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n19899)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16447_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(PWMdut_m3[9]), .B(PWMdut_m3[3]), .C(PWMdut_m3[4]), 
         .D(n11551), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_adj_149 (.A(PWMdut_m3[6]), .B(PWMdut_m3[7]), .Z(n10_adj_2389)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut_adj_149.init = 16'heeee;
    LUT4 i2_3_lut (.A(PWMdut_m3[2]), .B(PWMdut_m3[1]), .C(PWMdut_m3[0]), 
         .Z(n11551)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut.init = 16'hfefe;
    CCU2D cnt_2129_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18396), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2129_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2129_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2129_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2129_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18395), 
          .COUT(n18396), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2129_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2129_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2129_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2129_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18394), 
          .COUT(n18395), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2129_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2129_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2129_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2129_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18393), 
          .COUT(n18394), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2129_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2129_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2129_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2129_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18392), 
          .COUT(n18393), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2129_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2129_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2129_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2129_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18392), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2129_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2129_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2129_add_4_1.INJECT1_1 = "NO";
    LUT4 i7_4_lut_rep_333 (.A(PWMdut_m3[5]), .B(n14), .C(n10_adj_2389), 
         .D(PWMdut_m3[8]), .Z(n21434)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i7_4_lut_rep_333.init = 16'hfffe;
    LUT4 DutyCycle_9__I_0_i20_1_lut_4_lut (.A(PWMdut_m3[5]), .B(n14), .C(n10_adj_2389), 
         .D(PWMdut_m3[8]), .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam DutyCycle_9__I_0_i20_1_lut_4_lut.init = 16'h0001;
    FD1S3IX cnt_2129__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14214), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i0.GSR = "ENABLED";
    FD1S3IX cnt_2129__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14214), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i1.GSR = "ENABLED";
    FD1S3IX cnt_2129__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14214), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i2.GSR = "ENABLED";
    FD1S3IX cnt_2129__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14214), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i3.GSR = "ENABLED";
    FD1S3IX cnt_2129__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14214), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i4.GSR = "ENABLED";
    FD1S3IX cnt_2129__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14214), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i5.GSR = "ENABLED";
    FD1S3IX cnt_2129__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14214), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i6.GSR = "ENABLED";
    FD1S3IX cnt_2129__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14214), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i7.GSR = "ENABLED";
    FD1S3IX cnt_2129__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14214), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i8.GSR = "ENABLED";
    FD1S3IX cnt_2129__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14214), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2129__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR_U2
//

module PWMGENERATOR_U2 (PWMdut_m1, GND_net, PWM_m1, pwm_clk, LED1_c, 
            clkout_c_enable_362);
    input [9:0]PWMdut_m1;
    input GND_net;
    output PWM_m1;
    input pwm_clk;
    output LED1_c;
    input clkout_c_enable_362;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    
    wire n18346, n21433;
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    wire [9:0]n1;
    
    wire n18347, n18345, n7, n18344, n10, PWM_N_2176, n7_adj_2386, 
        n8, n11547, n18406;
    wire [9:0]n45;
    
    wire free_N_2188, n18405, n18404, n3853, n19903, n6, n14216, 
        n19869, n18403, n18402, n14, n18348;
    
    CCU2D sub_1802_add_2_7 (.A0(PWMdut_m1[5]), .B0(n21433), .C0(cnt[5]), 
          .D0(GND_net), .A1(n1[6]), .B1(n21433), .C1(cnt[6]), .D1(GND_net), 
          .CIN(n18346), .COUT(n18347));
    defparam sub_1802_add_2_7.INIT0 = 16'h8787;
    defparam sub_1802_add_2_7.INIT1 = 16'h8787;
    defparam sub_1802_add_2_7.INJECT1_0 = "NO";
    defparam sub_1802_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_5 (.A0(n1[3]), .B0(n21433), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(n21433), .C1(n7), .D1(PWMdut_m1[4]), .CIN(n18345), 
          .COUT(n18346));
    defparam sub_1802_add_2_5.INIT0 = 16'h8787;
    defparam sub_1802_add_2_5.INIT1 = 16'h5955;
    defparam sub_1802_add_2_5.INJECT1_0 = "NO";
    defparam sub_1802_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_3 (.A0(cnt[1]), .B0(n21433), .C0(n7), .D0(PWMdut_m1[1]), 
          .A1(cnt[2]), .B1(n21433), .C1(n7), .D1(PWMdut_m1[2]), .CIN(n18344), 
          .COUT(n18345));
    defparam sub_1802_add_2_3.INIT0 = 16'h5955;
    defparam sub_1802_add_2_3.INIT1 = 16'h5955;
    defparam sub_1802_add_2_3.INJECT1_0 = "NO";
    defparam sub_1802_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(n21433), .C1(n7), .D1(PWMdut_m1[0]), 
          .COUT(n18344));
    defparam sub_1802_add_2_1.INIT0 = 16'h0000;
    defparam sub_1802_add_2_1.INIT1 = 16'h5955;
    defparam sub_1802_add_2_1.INJECT1_0 = "NO";
    defparam sub_1802_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(PWMdut_m1[6]), .B(PWMdut_m1[7]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    FD1S3AX PWM_22 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m1)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=328, LSE_RLINE=328 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam PWM_22.GSR = "ENABLED";
    LUT4 i13267_2_lut (.A(PWMdut_m1[6]), .B(n7), .Z(n1[6])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13267_2_lut.init = 16'heeee;
    LUT4 i5_4_lut (.A(PWMdut_m1[9]), .B(n7_adj_2386), .C(PWMdut_m1[7]), 
         .D(n8), .Z(n7)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(PWMdut_m1[6]), .B(n11547), .C(PWMdut_m1[4]), .D(PWMdut_m1[3]), 
         .Z(n7_adj_2386)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut.init = 16'ha8a0;
    LUT4 i2_2_lut_adj_148 (.A(PWMdut_m1[5]), .B(PWMdut_m1[8]), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_148.init = 16'h8888;
    LUT4 i2_3_lut (.A(PWMdut_m1[2]), .B(PWMdut_m1[1]), .C(PWMdut_m1[0]), 
         .Z(n11547)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i13265_2_lut (.A(PWMdut_m1[3]), .B(n7), .Z(n1[3])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13265_2_lut.init = 16'heeee;
    CCU2D cnt_2127_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18406), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2127_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2127_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2127_add_4_11.INJECT1_1 = "NO";
    FD1P3AX free_21 (.D(free_N_2188), .SP(clkout_c_enable_362), .CK(pwm_clk), 
            .Q(LED1_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam free_21.GSR = "DISABLED";
    CCU2D cnt_2127_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18405), 
          .COUT(n18406), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2127_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2127_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2127_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2127_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18404), 
          .COUT(n18405), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2127_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2127_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2127_add_4_7.INJECT1_1 = "NO";
    LUT4 i1804_1_lut (.A(n3853), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1804_1_lut.init = 16'h5555;
    LUT4 i17198_4_lut (.A(cnt[2]), .B(n19903), .C(cnt[1]), .D(n6), .Z(n14216)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(77[6:16])
    defparam i17198_4_lut.init = 16'h0004;
    LUT4 i16451_3_lut (.A(cnt[6]), .B(n19869), .C(cnt[8]), .Z(n19903)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16451_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(cnt[4]), .B(cnt[0]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i16417_4_lut (.A(cnt[7]), .B(cnt[5]), .C(cnt[9]), .D(cnt[3]), 
         .Z(n19869)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16417_4_lut.init = 16'h8000;
    CCU2D cnt_2127_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18403), 
          .COUT(n18404), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2127_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2127_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2127_add_4_5.INJECT1_1 = "NO";
    LUT4 i13269_2_lut (.A(PWMdut_m1[8]), .B(n7), .Z(n1[8])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13269_2_lut.init = 16'heeee;
    CCU2D cnt_2127_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18402), 
          .COUT(n18403), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2127_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2127_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2127_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2127_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18402), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2127_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2127_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2127_add_4_1.INJECT1_1 = "NO";
    LUT4 i6_4_lut (.A(PWMdut_m1[9]), .B(PWMdut_m1[3]), .C(PWMdut_m1[4]), 
         .D(n11547), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut_rep_332 (.A(PWMdut_m1[5]), .B(n14), .C(n10), .D(PWMdut_m1[8]), 
         .Z(n21433)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i7_4_lut_rep_332.init = 16'hfffe;
    LUT4 DutyCycle_9__I_0_i20_1_lut_4_lut (.A(PWMdut_m1[5]), .B(n14), .C(n10), 
         .D(PWMdut_m1[8]), .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam DutyCycle_9__I_0_i20_1_lut_4_lut.init = 16'h0001;
    FD1S3IX cnt_2127__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14216), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i0.GSR = "ENABLED";
    FD1S3IX cnt_2127__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14216), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i1.GSR = "ENABLED";
    CCU2D sub_1802_add_2_11 (.A0(PWMdut_m1[9]), .B0(n21433), .C0(cnt[9]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18348), .S1(n3853));
    defparam sub_1802_add_2_11.INIT0 = 16'h8787;
    defparam sub_1802_add_2_11.INIT1 = 16'h0000;
    defparam sub_1802_add_2_11.INJECT1_0 = "NO";
    defparam sub_1802_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1802_add_2_9 (.A0(PWMdut_m1[7]), .B0(n21433), .C0(cnt[7]), 
          .D0(GND_net), .A1(n1[8]), .B1(n21433), .C1(cnt[8]), .D1(GND_net), 
          .CIN(n18347), .COUT(n18348));
    defparam sub_1802_add_2_9.INIT0 = 16'h8787;
    defparam sub_1802_add_2_9.INIT1 = 16'h8787;
    defparam sub_1802_add_2_9.INJECT1_0 = "NO";
    defparam sub_1802_add_2_9.INJECT1_1 = "NO";
    FD1S3IX cnt_2127__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14216), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i2.GSR = "ENABLED";
    FD1S3IX cnt_2127__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14216), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i3.GSR = "ENABLED";
    FD1S3IX cnt_2127__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14216), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i4.GSR = "ENABLED";
    FD1S3IX cnt_2127__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14216), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i5.GSR = "ENABLED";
    FD1S3IX cnt_2127__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14216), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i6.GSR = "ENABLED";
    FD1S3IX cnt_2127__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14216), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i7.GSR = "ENABLED";
    FD1S3IX cnt_2127__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14216), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i8.GSR = "ENABLED";
    FD1S3IX cnt_2127__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14216), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2127__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \PID(16000000,160000000,10000000) 
//

module \PID(16000000,160000000,10000000)  (speed_set_m2, GND_net, clk_N_875, 
            speed_set_m3, \subOut_24__N_1369[0] , speed_set_m1, speed_set_m4, 
            dir_m2, dir_m3, dir_m1, dir_m4, \speed_avg_m3[12] , \speed_avg_m2[12] , 
            \speed_avg_m1[12] , \speed_avg_m1[9] , \speed_avg_m1[8] , 
            \speed_avg_m1[7] , \speed_avg_m1[3] , \speed_avg_m1[19] , 
            \speed_avg_m2[19] , VCC_net, \speed_avg_m1[18] , \speed_avg_m2[18] , 
            \speed_avg_m1[17] , \speed_avg_m2[17] , \speed_avg_m1[16] , 
            \speed_avg_m2[16] , \speed_avg_m1[15] , \speed_avg_m2[15] , 
            \speed_avg_m1[14] , \speed_avg_m2[14] , \speed_avg_m1[13] , 
            \speed_avg_m2[13] , \speed_avg_m1[11] , \speed_avg_m2[11] , 
            \speed_avg_m1[10] , \speed_avg_m2[10] , \speed_avg_m1[6] , 
            \speed_avg_m2[6] , \speed_avg_m1[5] , \speed_avg_m2[5] , \speed_avg_m1[4] , 
            \speed_avg_m2[4] , \speed_avg_m1[2] , \speed_avg_m2[2] , \speed_avg_m3[9] , 
            \speed_avg_m2[9] , \speed_avg_m1[1] , \speed_avg_m2[1] , \speed_avg_m1[0] , 
            \speed_avg_m2[0] , n19649, \speed_avg_m3[8] , \speed_avg_m2[8] , 
            \speed_avg_m3[7] , \speed_avg_m2[7] , \speed_avg_m3[3] , \speed_avg_m2[3] , 
            \speed_avg_m4[19] , \speed_avg_m3[19] , \speed_avg_m4[18] , 
            \speed_avg_m3[18] , \speed_avg_m4[17] , \speed_avg_m3[17] , 
            \speed_avg_m4[16] , \speed_avg_m3[16] , \speed_avg_m4[15] , 
            \speed_avg_m3[15] , \speed_avg_m4[14] , \speed_avg_m3[14] , 
            \speed_avg_m4[13] , \speed_avg_m3[13] , \speed_avg_m4[11] , 
            \speed_avg_m3[11] , \speed_avg_m4[10] , \speed_avg_m3[10] , 
            \subOut_24__N_1369[1] , \subOut_24__N_1369[2] , \subOut_24__N_1369[3] , 
            \subOut_24__N_1369[4] , \subOut_24__N_1369[5] , \subOut_24__N_1369[6] , 
            \subOut_24__N_1369[7] , \subOut_24__N_1369[8] , \subOut_24__N_1369[9] , 
            \subOut_24__N_1369[10] , \subOut_24__N_1369[11] , \subOut_24__N_1369[12] , 
            \subOut_24__N_1369[13] , \subOut_24__N_1369[14] , \subOut_24__N_1369[15] , 
            \subOut_24__N_1369[16] , \subOut_24__N_1369[17] , \subOut_24__N_1369[18] , 
            \subOut_24__N_1369[19] , \subOut_24__N_1369[20] , \subOut_24__N_1369[21] , 
            \subOut_24__N_1369[24] , \speed_avg_m4[6] , \speed_avg_m3[6] , 
            \speed_avg_m4[5] , \speed_avg_m3[5] , \speed_avg_m4[4] , \speed_avg_m3[4] , 
            \speed_avg_m4[2] , \speed_avg_m3[2] , \speed_avg_m4[1] , \speed_avg_m3[1] , 
            \speed_avg_m4[0] , \speed_avg_m3[0] , \speed_avg_m4[12] , 
            \speed_avg_m4[9] , \speed_avg_m4[8] , \speed_avg_m4[7] , \speed_avg_m4[3] , 
            n22211, PWMdut_m4, PWMdut_m3, PWMdut_m2, PWMdut_m1, n4510, 
            n4512, n4511, n4514, n4513, n4516, n4515, n4518, n4517, 
            n4520, n4519, n4522, n4521, n4524, n4523, n4526, n4525, 
            n4528, n4527, n4530, n4529, n4531, n4485, n4484, n4487, 
            n4486, n4489, n4488, n4491, n4490, n4493, n4492, n4495, 
            n4494, n4497, n4496, n4499, n4498, n4501, n4500, n4503, 
            n4502, n4505, n4504, n4506);
    input [20:0]speed_set_m2;
    input GND_net;
    input clk_N_875;
    input [20:0]speed_set_m3;
    input \subOut_24__N_1369[0] ;
    input [20:0]speed_set_m1;
    input [20:0]speed_set_m4;
    output dir_m2;
    output dir_m3;
    output dir_m1;
    output dir_m4;
    input \speed_avg_m3[12] ;
    input \speed_avg_m2[12] ;
    input \speed_avg_m1[12] ;
    input \speed_avg_m1[9] ;
    input \speed_avg_m1[8] ;
    input \speed_avg_m1[7] ;
    input \speed_avg_m1[3] ;
    input \speed_avg_m1[19] ;
    input \speed_avg_m2[19] ;
    input VCC_net;
    input \speed_avg_m1[18] ;
    input \speed_avg_m2[18] ;
    input \speed_avg_m1[17] ;
    input \speed_avg_m2[17] ;
    input \speed_avg_m1[16] ;
    input \speed_avg_m2[16] ;
    input \speed_avg_m1[15] ;
    input \speed_avg_m2[15] ;
    input \speed_avg_m1[14] ;
    input \speed_avg_m2[14] ;
    input \speed_avg_m1[13] ;
    input \speed_avg_m2[13] ;
    input \speed_avg_m1[11] ;
    input \speed_avg_m2[11] ;
    input \speed_avg_m1[10] ;
    input \speed_avg_m2[10] ;
    input \speed_avg_m1[6] ;
    input \speed_avg_m2[6] ;
    input \speed_avg_m1[5] ;
    input \speed_avg_m2[5] ;
    input \speed_avg_m1[4] ;
    input \speed_avg_m2[4] ;
    input \speed_avg_m1[2] ;
    input \speed_avg_m2[2] ;
    input \speed_avg_m3[9] ;
    input \speed_avg_m2[9] ;
    input \speed_avg_m1[1] ;
    input \speed_avg_m2[1] ;
    input \speed_avg_m1[0] ;
    input \speed_avg_m2[0] ;
    output n19649;
    input \speed_avg_m3[8] ;
    input \speed_avg_m2[8] ;
    input \speed_avg_m3[7] ;
    input \speed_avg_m2[7] ;
    input \speed_avg_m3[3] ;
    input \speed_avg_m2[3] ;
    input \speed_avg_m4[19] ;
    input \speed_avg_m3[19] ;
    input \speed_avg_m4[18] ;
    input \speed_avg_m3[18] ;
    input \speed_avg_m4[17] ;
    input \speed_avg_m3[17] ;
    input \speed_avg_m4[16] ;
    input \speed_avg_m3[16] ;
    input \speed_avg_m4[15] ;
    input \speed_avg_m3[15] ;
    input \speed_avg_m4[14] ;
    input \speed_avg_m3[14] ;
    input \speed_avg_m4[13] ;
    input \speed_avg_m3[13] ;
    input \speed_avg_m4[11] ;
    input \speed_avg_m3[11] ;
    input \speed_avg_m4[10] ;
    input \speed_avg_m3[10] ;
    input \subOut_24__N_1369[1] ;
    input \subOut_24__N_1369[2] ;
    input \subOut_24__N_1369[3] ;
    input \subOut_24__N_1369[4] ;
    input \subOut_24__N_1369[5] ;
    input \subOut_24__N_1369[6] ;
    input \subOut_24__N_1369[7] ;
    input \subOut_24__N_1369[8] ;
    input \subOut_24__N_1369[9] ;
    input \subOut_24__N_1369[10] ;
    input \subOut_24__N_1369[11] ;
    input \subOut_24__N_1369[12] ;
    input \subOut_24__N_1369[13] ;
    input \subOut_24__N_1369[14] ;
    input \subOut_24__N_1369[15] ;
    input \subOut_24__N_1369[16] ;
    input \subOut_24__N_1369[17] ;
    input \subOut_24__N_1369[18] ;
    input \subOut_24__N_1369[19] ;
    input \subOut_24__N_1369[20] ;
    input \subOut_24__N_1369[21] ;
    input \subOut_24__N_1369[24] ;
    input \speed_avg_m4[6] ;
    input \speed_avg_m3[6] ;
    input \speed_avg_m4[5] ;
    input \speed_avg_m3[5] ;
    input \speed_avg_m4[4] ;
    input \speed_avg_m3[4] ;
    input \speed_avg_m4[2] ;
    input \speed_avg_m3[2] ;
    input \speed_avg_m4[1] ;
    input \speed_avg_m3[1] ;
    input \speed_avg_m4[0] ;
    input \speed_avg_m3[0] ;
    input \speed_avg_m4[12] ;
    input \speed_avg_m4[9] ;
    input \speed_avg_m4[8] ;
    input \speed_avg_m4[7] ;
    input \speed_avg_m4[3] ;
    input n22211;
    output [9:0]PWMdut_m4;
    output [9:0]PWMdut_m3;
    output [9:0]PWMdut_m2;
    output [9:0]PWMdut_m1;
    output n4510;
    output n4512;
    output n4511;
    output n4514;
    output n4513;
    output n4516;
    output n4515;
    output n4518;
    output n4517;
    output n4520;
    output n4519;
    output n4522;
    output n4521;
    output n4524;
    output n4523;
    output n4526;
    output n4525;
    output n4528;
    output n4527;
    output n4530;
    output n4529;
    output n4531;
    output n4485;
    output n4484;
    output n4487;
    output n4486;
    output n4489;
    output n4488;
    output n4491;
    output n4490;
    output n4493;
    output n4492;
    output n4495;
    output n4494;
    output n4497;
    output n4496;
    output n4499;
    output n4498;
    output n4501;
    output n4500;
    output n4503;
    output n4502;
    output n4505;
    output n4504;
    output n4506;
    
    wire clk_N_875 /* synthesis is_inv_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(30[4:14])
    wire [4:0]ss;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(96[9:11])
    
    wire n21492;
    wire [15:0]n1322;
    
    wire n8, n4, n10, n18534, n3656, n18533, n21471, n9, n21418, 
        n18413;
    wire [28:0]multOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(88[9:16])
    
    wire n16420;
    wire [28:0]addOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(92[9:15])
    wire [28:0]addIn2_28__N_1441;
    wire [28:0]n121;
    
    wire n18414, n18234, n5447, n5449;
    wire [21:0]n2373;
    
    wire n18235, n20118, n18532, n18531, n18412;
    wire [28:0]backOut0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(77[9:17])
    
    wire clk_N_875_enable_69;
    wire [28:0]Out3_28__N_1174;
    
    wire n22216, n21431, n21490, n22209, n21463, n16496, n42, 
        n5377, n22203, n18530;
    wire [28:0]backOut1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(78[9:17])
    
    wire clk_N_875_enable_41, n21498, n21505, n21504, n18529, n18471, 
        n5365, n21508, n21507, n18528, n21493, n21462, n21458, 
        clk_N_875_enable_392, n14360, clk_N_875_enable_303, n14388;
    wire [53:0]multOut_28__N_1412;
    
    wire n18527, n18526, n1068, n18470, n18469, n18525, n18411, 
        n18468, n18524, n5357, n5379, n18226;
    wire [15:0]n1301;
    wire [9:0]n2281;
    
    wire n18227, n18467, n18523, n15, n21494;
    wire [9:0]n2293;
    
    wire n30, n19107, n18522, n5375, n19101, n18410, n21407, n21406, 
        n21410, subIn1_24__N_1342, n11585, n3840;
    wire [28:0]intgOut0_28__N_1629;
    
    wire n18409;
    wire [28:0]Out0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(72[9:13])
    
    wire clk_N_875_enable_97;
    wire [28:0]Out1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(73[9:13])
    
    wire clk_N_875_enable_125;
    wire [28:0]Out2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(74[9:13])
    
    wire clk_N_875_enable_153;
    wire [28:0]Out3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(75[9:13])
    
    wire clk_N_875_enable_181;
    wire [28:0]backOut2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(79[9:17])
    
    wire clk_N_875_enable_209, n14;
    wire [28:0]backOut3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(80[9:17])
    
    wire clk_N_875_enable_237;
    wire [24:0]subOut;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(84[9:15])
    
    wire n18521, n5349, n5367, n18408, n18466, n18520, n18465, 
        n5359, n5351, n18464, n21464, n21467, n18519, n6, n21495, 
        n9_adj_2327, n18407;
    wire [9:0]n1458;
    
    wire n35, n21403, n19679, n18518, n18338;
    wire [15:0]n1364;
    wire [9:0]n2317;
    
    wire n18337, n18233, n5443, n5445, n18517, n5415, n21474, 
        n11644;
    wire [28:0]intgOut3;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(70[9:17])
    
    wire n14382, clk_N_875_enable_391, n14419, n21473;
    wire [28:0]n588;
    
    wire n5403, n21466, n49, n15773, n16542, n21499, n21470, n18225, 
        n18463, n18224, n18516, n18462, n5413, n9_adj_2328;
    wire [9:0]n1414;
    
    wire n18223, n18222, n9_adj_2329, n8_adj_2330, n18461, n10_adj_2331, 
        n18221, n8_adj_2332, n4_adj_2333, n18220, n18215, n18216;
    wire [28:0]intgOut0;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(67[9:17])
    wire [28:0]n648;
    wire [28:0]n678;
    
    wire n18217, n18218, n19674, n18219, n5884, n14410, subIn1_24__N_1534, 
        dirout_m3_N_1949, subIn1_24__N_1347, dirout_m4_N_1952;
    wire [28:0]backOut2_28__N_1845;
    
    wire n18460;
    wire [28:0]Out0_28__N_1087;
    wire [28:0]Out2_28__N_1145;
    
    wire n18273;
    wire [28:0]backOut3_28__N_1874;
    
    wire n5556, n22204;
    wire [20:0]subIn2_24__N_1535;
    
    wire n16258, n19662, n21424, n5868;
    wire [20:0]subIn2_24__N_1348;
    wire [23:0]multIn2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(87[9:16])
    
    wire mult_29s_25s_0_pp_1_2, mult_29s_25s_0_pp_2_4, mult_29s_25s_0_pp_3_6, 
        mult_29s_25s_0_pp_4_8, mult_29s_25s_0_pp_5_10, mult_29s_25s_0_pp_6_12, 
        mult_29s_25s_0_pp_7_14, mult_29s_25s_0_pp_8_16, mult_29s_25s_0_pp_9_18, 
        mult_29s_25s_0_pp_10_20, mult_29s_25s_0_pp_11_22, mult_29s_25s_0_pp_12_24, 
        mult_29s_25s_0_pp_12_25, mult_29s_25s_0_pp_12_26, mult_29s_25s_0_pp_12_27, 
        mult_29s_25s_0_pp_12_28, mult_29s_25s_0_cin_lr_2, mult_29s_25s_0_cin_lr_4, 
        mult_29s_25s_0_cin_lr_6, mult_29s_25s_0_cin_lr_8, mult_29s_25s_0_cin_lr_10, 
        mult_29s_25s_0_cin_lr_12, mult_29s_25s_0_cin_lr_14, mult_29s_25s_0_cin_lr_16, 
        mult_29s_25s_0_cin_lr_18, mult_29s_25s_0_cin_lr_20, mult_29s_25s_0_cin_lr_22, 
        co_mult_29s_25s_0_0_1, mult_29s_25s_0_pp_0_2, co_mult_29s_25s_0_0_2, 
        s_mult_29s_25s_0_0_4, mult_29s_25s_0_pp_0_4, mult_29s_25s_0_pp_0_3, 
        mult_29s_25s_0_pp_1_4, mult_29s_25s_0_pp_1_3, co_mult_29s_25s_0_0_3, 
        s_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_6, mult_29s_25s_0_pp_0_6, 
        mult_29s_25s_0_pp_0_5, mult_29s_25s_0_pp_1_6, mult_29s_25s_0_pp_1_5, 
        co_mult_29s_25s_0_0_4, s_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_8, 
        mult_29s_25s_0_pp_0_8, mult_29s_25s_0_pp_0_7, mult_29s_25s_0_pp_1_8, 
        mult_29s_25s_0_pp_1_7, co_mult_29s_25s_0_0_5, s_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_10, mult_29s_25s_0_pp_0_10, mult_29s_25s_0_pp_0_9, 
        mult_29s_25s_0_pp_1_10, mult_29s_25s_0_pp_1_9, co_mult_29s_25s_0_0_6, 
        s_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_12, mult_29s_25s_0_pp_0_12, 
        mult_29s_25s_0_pp_0_11, mult_29s_25s_0_pp_1_12, mult_29s_25s_0_pp_1_11, 
        co_mult_29s_25s_0_0_7, s_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_14, 
        mult_29s_25s_0_pp_0_14, mult_29s_25s_0_pp_0_13, mult_29s_25s_0_pp_1_14, 
        mult_29s_25s_0_pp_1_13, co_mult_29s_25s_0_0_8, s_mult_29s_25s_0_0_15, 
        s_mult_29s_25s_0_0_16, mult_29s_25s_0_pp_0_16, mult_29s_25s_0_pp_0_15, 
        mult_29s_25s_0_pp_1_16, mult_29s_25s_0_pp_1_15, co_mult_29s_25s_0_0_9, 
        s_mult_29s_25s_0_0_17, s_mult_29s_25s_0_0_18, mult_29s_25s_0_pp_0_18, 
        mult_29s_25s_0_pp_0_17, mult_29s_25s_0_pp_1_18, mult_29s_25s_0_pp_1_17, 
        co_mult_29s_25s_0_0_10, s_mult_29s_25s_0_0_19, s_mult_29s_25s_0_0_20, 
        mult_29s_25s_0_pp_0_20, mult_29s_25s_0_pp_0_19, mult_29s_25s_0_pp_1_20, 
        mult_29s_25s_0_pp_1_19, co_mult_29s_25s_0_0_11, s_mult_29s_25s_0_0_21, 
        s_mult_29s_25s_0_0_22, mult_29s_25s_0_pp_0_22, mult_29s_25s_0_pp_0_21, 
        mult_29s_25s_0_pp_1_22, mult_29s_25s_0_pp_1_21, co_mult_29s_25s_0_0_12, 
        s_mult_29s_25s_0_0_23, s_mult_29s_25s_0_0_24, mult_29s_25s_0_pp_0_24, 
        mult_29s_25s_0_pp_0_23, mult_29s_25s_0_pp_1_24, mult_29s_25s_0_pp_1_23, 
        co_mult_29s_25s_0_0_13, s_mult_29s_25s_0_0_25, s_mult_29s_25s_0_0_26, 
        mult_29s_25s_0_pp_0_26, mult_29s_25s_0_pp_0_25, mult_29s_25s_0_pp_1_26, 
        mult_29s_25s_0_pp_1_25, s_mult_29s_25s_0_0_27, s_mult_29s_25s_0_0_28, 
        mult_29s_25s_0_pp_0_28, mult_29s_25s_0_pp_0_27, mult_29s_25s_0_pp_1_28, 
        mult_29s_25s_0_pp_1_27, co_mult_29s_25s_0_1_1, s_mult_29s_25s_0_1_6, 
        mult_29s_25s_0_pp_2_6, co_mult_29s_25s_0_1_2, s_mult_29s_25s_0_1_7, 
        s_mult_29s_25s_0_1_8, mult_29s_25s_0_pp_2_8, mult_29s_25s_0_pp_2_7, 
        mult_29s_25s_0_pp_3_8, mult_29s_25s_0_pp_3_7, co_mult_29s_25s_0_1_3, 
        s_mult_29s_25s_0_1_9, s_mult_29s_25s_0_1_10, mult_29s_25s_0_pp_2_10, 
        mult_29s_25s_0_pp_2_9, mult_29s_25s_0_pp_3_10, mult_29s_25s_0_pp_3_9, 
        co_mult_29s_25s_0_1_4, s_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_12, 
        mult_29s_25s_0_pp_2_12, mult_29s_25s_0_pp_2_11, mult_29s_25s_0_pp_3_12, 
        mult_29s_25s_0_pp_3_11, co_mult_29s_25s_0_1_5, s_mult_29s_25s_0_1_13, 
        s_mult_29s_25s_0_1_14, mult_29s_25s_0_pp_2_14, mult_29s_25s_0_pp_2_13, 
        mult_29s_25s_0_pp_3_14, mult_29s_25s_0_pp_3_13, co_mult_29s_25s_0_1_6, 
        s_mult_29s_25s_0_1_15, s_mult_29s_25s_0_1_16, mult_29s_25s_0_pp_2_16, 
        mult_29s_25s_0_pp_2_15, mult_29s_25s_0_pp_3_16, mult_29s_25s_0_pp_3_15, 
        co_mult_29s_25s_0_1_7, s_mult_29s_25s_0_1_17, s_mult_29s_25s_0_1_18, 
        mult_29s_25s_0_pp_2_18, mult_29s_25s_0_pp_2_17, mult_29s_25s_0_pp_3_18, 
        mult_29s_25s_0_pp_3_17, co_mult_29s_25s_0_1_8, s_mult_29s_25s_0_1_19, 
        s_mult_29s_25s_0_1_20, mult_29s_25s_0_pp_2_20, mult_29s_25s_0_pp_2_19, 
        mult_29s_25s_0_pp_3_20, mult_29s_25s_0_pp_3_19, co_mult_29s_25s_0_1_9, 
        s_mult_29s_25s_0_1_21, s_mult_29s_25s_0_1_22, mult_29s_25s_0_pp_2_22, 
        mult_29s_25s_0_pp_2_21, mult_29s_25s_0_pp_3_22, mult_29s_25s_0_pp_3_21, 
        co_mult_29s_25s_0_1_10, s_mult_29s_25s_0_1_23, s_mult_29s_25s_0_1_24, 
        mult_29s_25s_0_pp_2_24, mult_29s_25s_0_pp_2_23, mult_29s_25s_0_pp_3_24, 
        mult_29s_25s_0_pp_3_23, co_mult_29s_25s_0_1_11, s_mult_29s_25s_0_1_25, 
        s_mult_29s_25s_0_1_26, mult_29s_25s_0_pp_2_26, mult_29s_25s_0_pp_2_25, 
        mult_29s_25s_0_pp_3_26, mult_29s_25s_0_pp_3_25, s_mult_29s_25s_0_1_27, 
        s_mult_29s_25s_0_1_28, mult_29s_25s_0_pp_2_28, mult_29s_25s_0_pp_2_27, 
        mult_29s_25s_0_pp_3_28, mult_29s_25s_0_pp_3_27, co_mult_29s_25s_0_2_1, 
        s_mult_29s_25s_0_2_10, mult_29s_25s_0_pp_4_10, co_mult_29s_25s_0_2_2, 
        s_mult_29s_25s_0_2_12, s_mult_29s_25s_0_2_11, mult_29s_25s_0_pp_4_12, 
        mult_29s_25s_0_pp_4_11, mult_29s_25s_0_pp_5_12, mult_29s_25s_0_pp_5_11, 
        co_mult_29s_25s_0_2_3, s_mult_29s_25s_0_2_13, s_mult_29s_25s_0_2_14, 
        mult_29s_25s_0_pp_4_14, mult_29s_25s_0_pp_4_13, mult_29s_25s_0_pp_5_14, 
        mult_29s_25s_0_pp_5_13, co_mult_29s_25s_0_2_4, s_mult_29s_25s_0_2_15, 
        s_mult_29s_25s_0_2_16, mult_29s_25s_0_pp_4_16, mult_29s_25s_0_pp_4_15, 
        mult_29s_25s_0_pp_5_16, mult_29s_25s_0_pp_5_15, co_mult_29s_25s_0_2_5, 
        s_mult_29s_25s_0_2_17, s_mult_29s_25s_0_2_18, mult_29s_25s_0_pp_4_18, 
        mult_29s_25s_0_pp_4_17, mult_29s_25s_0_pp_5_18, mult_29s_25s_0_pp_5_17, 
        co_mult_29s_25s_0_2_6, s_mult_29s_25s_0_2_19, s_mult_29s_25s_0_2_20, 
        mult_29s_25s_0_pp_4_20, mult_29s_25s_0_pp_4_19, mult_29s_25s_0_pp_5_20, 
        mult_29s_25s_0_pp_5_19, co_mult_29s_25s_0_2_7, s_mult_29s_25s_0_2_21, 
        s_mult_29s_25s_0_2_22, mult_29s_25s_0_pp_4_22, mult_29s_25s_0_pp_4_21, 
        mult_29s_25s_0_pp_5_22, mult_29s_25s_0_pp_5_21, co_mult_29s_25s_0_2_8, 
        s_mult_29s_25s_0_2_23, s_mult_29s_25s_0_2_24, mult_29s_25s_0_pp_4_24, 
        mult_29s_25s_0_pp_4_23, mult_29s_25s_0_pp_5_24, mult_29s_25s_0_pp_5_23, 
        co_mult_29s_25s_0_2_9, s_mult_29s_25s_0_2_25, s_mult_29s_25s_0_2_26, 
        mult_29s_25s_0_pp_4_26, mult_29s_25s_0_pp_4_25, mult_29s_25s_0_pp_5_26, 
        mult_29s_25s_0_pp_5_25, s_mult_29s_25s_0_2_27, s_mult_29s_25s_0_2_28, 
        mult_29s_25s_0_pp_4_28, mult_29s_25s_0_pp_4_27, mult_29s_25s_0_pp_5_28, 
        mult_29s_25s_0_pp_5_27, co_mult_29s_25s_0_3_1, s_mult_29s_25s_0_3_14, 
        mult_29s_25s_0_pp_6_14, co_mult_29s_25s_0_3_2, s_mult_29s_25s_0_3_15, 
        s_mult_29s_25s_0_3_16, mult_29s_25s_0_pp_6_16, mult_29s_25s_0_pp_6_15, 
        mult_29s_25s_0_pp_7_16, mult_29s_25s_0_pp_7_15, co_mult_29s_25s_0_3_3, 
        s_mult_29s_25s_0_3_17, s_mult_29s_25s_0_3_18, mult_29s_25s_0_pp_6_18, 
        mult_29s_25s_0_pp_6_17, mult_29s_25s_0_pp_7_18, mult_29s_25s_0_pp_7_17, 
        co_mult_29s_25s_0_3_4, s_mult_29s_25s_0_3_19, s_mult_29s_25s_0_3_20, 
        mult_29s_25s_0_pp_6_20, mult_29s_25s_0_pp_6_19, mult_29s_25s_0_pp_7_20, 
        mult_29s_25s_0_pp_7_19, co_mult_29s_25s_0_3_5, s_mult_29s_25s_0_3_21, 
        s_mult_29s_25s_0_3_22, mult_29s_25s_0_pp_6_22, mult_29s_25s_0_pp_6_21, 
        mult_29s_25s_0_pp_7_22, mult_29s_25s_0_pp_7_21, co_mult_29s_25s_0_3_6, 
        s_mult_29s_25s_0_3_23, s_mult_29s_25s_0_3_24, mult_29s_25s_0_pp_6_24, 
        mult_29s_25s_0_pp_6_23, mult_29s_25s_0_pp_7_24, mult_29s_25s_0_pp_7_23, 
        co_mult_29s_25s_0_3_7, s_mult_29s_25s_0_3_25, s_mult_29s_25s_0_3_26, 
        mult_29s_25s_0_pp_6_26, mult_29s_25s_0_pp_6_25, mult_29s_25s_0_pp_7_26, 
        mult_29s_25s_0_pp_7_25, s_mult_29s_25s_0_3_27, s_mult_29s_25s_0_3_28, 
        mult_29s_25s_0_pp_6_28, mult_29s_25s_0_pp_6_27, mult_29s_25s_0_pp_7_28, 
        mult_29s_25s_0_pp_7_27, co_mult_29s_25s_0_4_1, s_mult_29s_25s_0_4_18, 
        mult_29s_25s_0_pp_8_18, co_mult_29s_25s_0_4_2, s_mult_29s_25s_0_4_20, 
        s_mult_29s_25s_0_4_19, mult_29s_25s_0_pp_8_20, mult_29s_25s_0_pp_8_19, 
        mult_29s_25s_0_pp_9_20, mult_29s_25s_0_pp_9_19, co_mult_29s_25s_0_4_3, 
        s_mult_29s_25s_0_4_21, s_mult_29s_25s_0_4_22, mult_29s_25s_0_pp_8_22, 
        mult_29s_25s_0_pp_8_21, mult_29s_25s_0_pp_9_22, mult_29s_25s_0_pp_9_21, 
        co_mult_29s_25s_0_4_4, s_mult_29s_25s_0_4_23, s_mult_29s_25s_0_4_24, 
        mult_29s_25s_0_pp_8_24, mult_29s_25s_0_pp_8_23, mult_29s_25s_0_pp_9_24, 
        mult_29s_25s_0_pp_9_23, co_mult_29s_25s_0_4_5, s_mult_29s_25s_0_4_25, 
        s_mult_29s_25s_0_4_26, mult_29s_25s_0_pp_8_26, mult_29s_25s_0_pp_8_25, 
        mult_29s_25s_0_pp_9_26, mult_29s_25s_0_pp_9_25, s_mult_29s_25s_0_4_27, 
        s_mult_29s_25s_0_4_28, mult_29s_25s_0_pp_8_28, mult_29s_25s_0_pp_8_27, 
        mult_29s_25s_0_pp_9_28, mult_29s_25s_0_pp_9_27, co_mult_29s_25s_0_5_1, 
        s_mult_29s_25s_0_5_22, mult_29s_25s_0_pp_10_22, co_mult_29s_25s_0_5_2, 
        s_mult_29s_25s_0_5_23, s_mult_29s_25s_0_5_24, mult_29s_25s_0_pp_10_24, 
        mult_29s_25s_0_pp_10_23, mult_29s_25s_0_pp_11_24, mult_29s_25s_0_pp_11_23, 
        co_mult_29s_25s_0_5_3, s_mult_29s_25s_0_5_25, s_mult_29s_25s_0_5_26, 
        mult_29s_25s_0_pp_10_26, mult_29s_25s_0_pp_10_25, mult_29s_25s_0_pp_11_26, 
        mult_29s_25s_0_pp_11_25, s_mult_29s_25s_0_5_27, s_mult_29s_25s_0_5_28, 
        mult_29s_25s_0_pp_10_28, mult_29s_25s_0_pp_10_27, mult_29s_25s_0_pp_11_28, 
        mult_29s_25s_0_pp_11_27, co_mult_29s_25s_0_6_1, s_mult_29s_25s_0_6_24, 
        co_mult_29s_25s_0_6_2, s_mult_29s_25s_0_6_25, s_mult_29s_25s_0_6_26, 
        s_mult_29s_25s_0_6_27, s_mult_29s_25s_0_6_28, co_mult_29s_25s_0_7_1, 
        co_mult_29s_25s_0_7_2, mult_29s_25s_0_pp_2_5, co_mult_29s_25s_0_7_3, 
        s_mult_29s_25s_0_7_8, co_mult_29s_25s_0_7_4, s_mult_29s_25s_0_7_9, 
        s_mult_29s_25s_0_7_10, co_mult_29s_25s_0_7_5, s_mult_29s_25s_0_7_11, 
        s_mult_29s_25s_0_7_12, co_mult_29s_25s_0_7_6, s_mult_29s_25s_0_7_13, 
        s_mult_29s_25s_0_7_14, co_mult_29s_25s_0_7_7, s_mult_29s_25s_0_7_15, 
        s_mult_29s_25s_0_7_16, co_mult_29s_25s_0_7_8, s_mult_29s_25s_0_7_17, 
        s_mult_29s_25s_0_7_18, co_mult_29s_25s_0_7_9, s_mult_29s_25s_0_7_19, 
        s_mult_29s_25s_0_7_20, co_mult_29s_25s_0_7_10, s_mult_29s_25s_0_7_21, 
        s_mult_29s_25s_0_7_22, co_mult_29s_25s_0_7_11, s_mult_29s_25s_0_7_23, 
        s_mult_29s_25s_0_7_24, co_mult_29s_25s_0_7_12, s_mult_29s_25s_0_7_25, 
        s_mult_29s_25s_0_7_26, s_mult_29s_25s_0_7_27, s_mult_29s_25s_0_7_28, 
        co_mult_29s_25s_0_8_1, s_mult_29s_25s_0_8_12, co_mult_29s_25s_0_8_2, 
        s_mult_29s_25s_0_8_13, s_mult_29s_25s_0_8_14, mult_29s_25s_0_pp_6_13, 
        co_mult_29s_25s_0_8_3, s_mult_29s_25s_0_8_15, s_mult_29s_25s_0_8_16, 
        co_mult_29s_25s_0_8_4, s_mult_29s_25s_0_8_17, s_mult_29s_25s_0_8_18, 
        co_mult_29s_25s_0_8_5, s_mult_29s_25s_0_8_19, s_mult_29s_25s_0_8_20, 
        co_mult_29s_25s_0_8_6, s_mult_29s_25s_0_8_21, s_mult_29s_25s_0_8_22, 
        co_mult_29s_25s_0_8_7, s_mult_29s_25s_0_8_23, s_mult_29s_25s_0_8_24, 
        co_mult_29s_25s_0_8_8, s_mult_29s_25s_0_8_25, s_mult_29s_25s_0_8_26, 
        s_mult_29s_25s_0_8_27, s_mult_29s_25s_0_8_28, co_mult_29s_25s_0_9_1, 
        s_mult_29s_25s_0_9_20, co_mult_29s_25s_0_9_2, s_mult_29s_25s_0_9_21, 
        s_mult_29s_25s_0_9_22, mult_29s_25s_0_pp_10_21, co_mult_29s_25s_0_9_3, 
        s_mult_29s_25s_0_9_24, s_mult_29s_25s_0_9_23, co_mult_29s_25s_0_9_4, 
        s_mult_29s_25s_0_9_25, s_mult_29s_25s_0_9_26, s_mult_29s_25s_0_9_27, 
        s_mult_29s_25s_0_9_28, co_mult_29s_25s_0_10_1, co_mult_29s_25s_0_10_2, 
        mult_29s_25s_0_pp_4_9, co_mult_29s_25s_0_10_3, co_mult_29s_25s_0_10_4, 
        co_mult_29s_25s_0_10_5, s_mult_29s_25s_0_10_16, co_mult_29s_25s_0_10_6, 
        s_mult_29s_25s_0_10_17, s_mult_29s_25s_0_10_18, co_mult_29s_25s_0_10_7, 
        s_mult_29s_25s_0_10_19, s_mult_29s_25s_0_10_20, co_mult_29s_25s_0_10_8, 
        s_mult_29s_25s_0_10_21, s_mult_29s_25s_0_10_22, co_mult_29s_25s_0_10_9, 
        s_mult_29s_25s_0_10_23, s_mult_29s_25s_0_10_24, co_mult_29s_25s_0_10_10, 
        s_mult_29s_25s_0_10_25, s_mult_29s_25s_0_10_26, s_mult_29s_25s_0_10_27, 
        s_mult_29s_25s_0_10_28, n18272, co_mult_29s_25s_0_11_1, s_mult_29s_25s_0_11_24, 
        co_mult_29s_25s_0_11_2, s_mult_29s_25s_0_11_25, s_mult_29s_25s_0_11_26, 
        s_mult_29s_25s_0_11_27, s_mult_29s_25s_0_11_28, n5870, co_t_mult_29s_25s_0_12_1, 
        co_t_mult_29s_25s_0_12_2, mult_29s_25s_0_pp_8_17, co_t_mult_29s_25s_0_12_3, 
        co_t_mult_29s_25s_0_12_4, co_t_mult_29s_25s_0_12_5, co_t_mult_29s_25s_0_12_6, 
        mult_29s_25s_0_cin_lr_0, mco, mco_1, mco_2, mco_3, mco_4, 
        mco_5, mco_6, mco_7, mco_8, mco_9, mco_10, mco_11, mco_12, 
        mco_14, mco_15, mco_16, mco_17, mco_18, mco_19, mco_20, 
        mco_21, mco_22, mco_23, mco_24, mco_25, mco_28, mco_29, 
        mco_30, mco_31, mco_32, mco_33, mco_34, mco_35, mco_36, 
        mco_37, mco_38, mco_42, mco_43, mco_44, mco_45, mco_46, 
        mco_47, mco_48, mco_49, mco_50, mco_51, mco_56, mco_57, 
        mco_58, mco_59, mco_60, mco_61, mco_62, mco_63, mco_64, 
        mco_70, mco_71, mco_72, mco_73, mco_74, mco_75, mco_76, 
        mco_77, mco_84, mco_85, mco_86, mco_87, mco_88, mco_89, 
        mco_90, mco_98, mco_99, mco_100, mco_101, mco_102, mco_103, 
        mco_112, mco_113, mco_114, mco_115, mco_116, mco_126, mco_127, 
        mco_128, mco_129, mco_140, mco_141, mco_142, mco_154, mco_155, 
        n5872, n21409, n15757, n21408, n56, n16223, n21427, n15143, 
        n21404, n21405, n5874, n21438, clk_N_875_enable_387, n14299, 
        n5876, n21448, n4389, n14_adj_2334, n10_adj_2335, n18754, 
        n6_adj_2336, n18755, n5878, n5880, n14_adj_2337, n10_adj_2338, 
        n18757, n6_adj_2339, n18758, n21440, clk_N_875_enable_359, 
        n15130, n5882, n16670, n16296, n3704, n35_adj_2340, n40, 
        n36, n4_adj_2341, n38, n32, n5886, n14_adj_2342, n10_adj_2343, 
        n18721, n34, n24, n6_adj_2344, n18722, n16678, n18698, 
        n5409, n35_adj_2345, n40_adj_2346, n36_adj_2347, n4_adj_2348, 
        n5419, n5423, n5421, n38_adj_2349, n32_adj_2350, n5888, 
        n34_adj_2351, n24_adj_2352, n5405, n5890, n16301, n19646, 
        n5393, n16674, n19672, n3608, n35_adj_2353, n40_adj_2354, 
        n36_adj_2355, n4_adj_2356, n38_adj_2357, n32_adj_2358, n21430;
    wire [28:0]n558;
    
    wire n5892, n34_adj_2359, n24_adj_2360, n3752, n35_adj_2361, n40_adj_2362, 
        n36_adj_2363, n4_adj_2364, n38_adj_2365, n32_adj_2366, n20157, 
        n34_adj_2367, n24_adj_2368, n5894, n14_adj_2369, n10_adj_2370, 
        n18759, n6_adj_2371, n18760, n5411, n21420;
    wire [20:0]n367;
    
    wire n5896, n21446, n21444, n21432, n20127, n5898, n5900, 
        n21475, n5902, n21491, n14304, n14332, n5904, n20388, 
        n5908, n21472, n5391, n21443, n5347, n18232, n5439, n5441, 
        n18271, n18270, n18231, n5435, n5437, n5399, n18459, n18458, 
        n18336, n18335, n18457, n18456, n5433, n14414, n18455, 
        n18334, n18454, n5369, n8_adj_2372, n21465, n3680, n18453, 
        n18452, n18451, n18450, n18449, n18448, n18447, n3632, 
        n18446, n18445, n18230, n18229;
    wire [15:0]n1343;
    wire [9:0]n2305;
    
    wire n9_adj_2373;
    wire [9:0]n1502;
    wire [28:0]intgOut1;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(68[9:17])
    wire [28:0]intgOut2;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(69[9:17])
    
    wire n18333, n18269, n18268, n18267, n18228, n18266, n18332, 
        n18331, n18330, n18329, n18444, n18265, n18264, n18263, 
        n18262, n18328, n18327, n18326, n18443, n18261, n18260;
    wire [21:0]n2613;
    
    wire n5407, n18259, n18258, n18325, n18324, n18442, n18257, 
        n18256, n18255, n18441, n18440, n18497, n18254, n18496, 
        n18439, n18253, n18252, n18251, n18250, n18438, n18495, 
        n18249, n18437, n18436, n18494, n5401, n5397, n3776, n18435, 
        n5361, n5395, n18434, n18433, n18493, n5417, n5427, n30_adj_2374, 
        n19131, n18248, n9_adj_2375, n7, n18492, n18491, n10_adj_2376, 
        n8_adj_2377, n4_adj_2378, n19125, n2565, n19119;
    wire [9:0]n1546;
    
    wire n5355, n5373, n5387, n5383, n5429, n5381, n5363, n5353, 
        n5371, n5473, n5385, n5471, n5425, n5469, n5467, n5465, 
        n14437, n5463, n5461, n5459, n5457, n18432, n18247, n5455, 
        n5453, n18246, n5451, n18431, n18430, n18490, n18245, 
        n18303, n18302, n9_adj_2379, n5345, n5557, n5869, n5871, 
        n5873, n5875, n18301, n18300, n18244, n5877, n5879, n5881, 
        n5883, n5885, n5887, n5889, n5891, n5893, n5895, n18299, 
        n18298, n18297, n18243, n5897, n5899, n5901, n9_adj_2380, 
        n8_adj_2381, n5903, n5905, n5909, n18296;
    wire [28:0]n618;
    wire [28:0]addIn2_28__N_1571;
    
    wire n10_adj_2382, n8_adj_2383, n4_adj_2384, n18489, n18488, n14428, 
        n19113, n20374, n4447, n4450, n4451, n18487, n4452, n4456, 
        n4440, n4441, n4442, n4443, n4444, n18295, n4445, n4446, 
        n4448, n4449, n4453, n4454, n4455, n4457, n4458, n4459, 
        n18294, n18486, n18485, n18484, n18242, n18483, n18241, 
        n18633, n18632, n18631, n18630, n18629, n18628, n18627, 
        n18626, n18625, n18482, n18481, n18480, n18624, n3728, 
        n18420, n18419, n18240, n18239, n18613, n18612, n18611, 
        n18610, n18609, n18608, n18607, n18606, n18605, n18604, 
        n18238, n18593, n18592, n18591, n18590, n18589, n18588, 
        n18587, n18586, n18585, n18584, n7_adj_2385, n18583, n18581, 
        n18580, n18579, n18578, n18577, n18576, n18575, n18574, 
        n18573, n18572, n18571, n18552, n18551, n18550, n18549, 
        n18548, n18547, n18546, n18545, n18544, n18543, n18542, 
        n18541, n18540, n18539, n18538, n18537, n18536, n18535, 
        n18237, n18418, n18417, n18416, n18236, n18415;
    
    LUT4 i1_2_lut_rep_391 (.A(ss[2]), .B(ss[1]), .Z(n21492)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_391.init = 16'heeee;
    LUT4 i4_4_lut (.A(n1322[6]), .B(n8), .C(n1322[4]), .D(n4), .Z(n10)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut.init = 16'hfeee;
    CCU2D add_15124_17 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18534), .S1(n3656));
    defparam add_15124_17.INIT0 = 16'h5555;
    defparam add_15124_17.INIT1 = 16'h0000;
    defparam add_15124_17.INJECT1_0 = "NO";
    defparam add_15124_17.INJECT1_1 = "NO";
    CCU2D add_15124_15 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18533), .COUT(n18534));
    defparam add_15124_15.INIT0 = 16'hf555;
    defparam add_15124_15.INIT1 = 16'hf555;
    defparam add_15124_15.INJECT1_0 = "NO";
    defparam add_15124_15.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_317_4_lut_4_lut_4_lut (.A(ss[1]), .B(n21471), .C(n9), 
         .Z(n21418)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(172[20:27])
    defparam i2_3_lut_rep_317_4_lut_4_lut_4_lut.init = 16'hd0d0;
    CCU2D addOut_2126_add_4_15 (.A0(multOut[13]), .B0(n16420), .C0(addOut[13]), 
          .D0(addIn2_28__N_1441[13]), .A1(multOut[14]), .B1(n16420), .C1(addOut[14]), 
          .D1(addIn2_28__N_1441[14]), .CIN(n18413), .COUT(n18414), .S0(n121[13]), 
          .S1(n121[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_15.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_15.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_15.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_15.INJECT1_1 = "NO";
    CCU2D add_1212_9 (.A0(n5447), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5449), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18234), 
          .COUT(n18235), .S0(n2373[7]), .S1(n2373[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_9.INIT0 = 16'hf555;
    defparam add_1212_9.INIT1 = 16'hf555;
    defparam add_1212_9.INJECT1_0 = "NO";
    defparam add_1212_9.INJECT1_1 = "NO";
    LUT4 i16652_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut (.A(ss[0]), .B(n21471), 
         .C(n9), .Z(n20118)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam i16652_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hd0d0;
    CCU2D add_15124_13 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18532), .COUT(n18533));
    defparam add_15124_13.INIT0 = 16'hf555;
    defparam add_15124_13.INIT1 = 16'hf555;
    defparam add_15124_13.INJECT1_0 = "NO";
    defparam add_15124_13.INJECT1_1 = "NO";
    CCU2D add_15124_11 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18531), .COUT(n18532));
    defparam add_15124_11.INIT0 = 16'hf555;
    defparam add_15124_11.INIT1 = 16'hf555;
    defparam add_15124_11.INJECT1_0 = "NO";
    defparam add_15124_11.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_13 (.A0(multOut[11]), .B0(n16420), .C0(addOut[11]), 
          .D0(addIn2_28__N_1441[11]), .A1(multOut[12]), .B1(n16420), .C1(addOut[12]), 
          .D1(addIn2_28__N_1441[12]), .CIN(n18412), .COUT(n18413), .S0(n121[11]), 
          .S1(n121[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_13.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_13.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_13.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_13.INJECT1_1 = "NO";
    FD1P3AX backOut0_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_330_3_lut_4_lut (.A(ss[2]), .B(ss[1]), .C(n22216), 
         .D(ss[3]), .Z(n21431)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C+!(D))))) */ ;
    defparam i1_2_lut_rep_330_3_lut_4_lut.init = 16'h010e;
    FD1S3IX ss_i0 (.D(n21490), .CK(clk_N_875), .CD(ss[4]), .Q(ss[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_362_3_lut_4_lut (.A(n22209), .B(ss[1]), .C(ss[3]), 
         .D(ss[0]), .Z(n21463)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_362_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1222_i16_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[15]), 
         .D(speed_set_m3[15]), .Z(n5377)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i16_3_lut_4_lut.init = 16'hfb40;
    FD1S3IX ss_i1 (.D(n22203), .CK(clk_N_875), .CD(ss[4]), .Q(ss[1]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i1.GSR = "ENABLED";
    CCU2D add_15124_9 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18530), .COUT(n18531));
    defparam add_15124_9.INIT0 = 16'hf555;
    defparam add_15124_9.INIT1 = 16'h0aaa;
    defparam add_15124_9.INJECT1_0 = "NO";
    defparam add_15124_9.INJECT1_1 = "NO";
    FD1P3AX backOut1_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i0.GSR = "DISABLED";
    LUT4 i1869_2_lut_rep_399 (.A(ss[0]), .B(ss[1]), .Z(n22203)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1869_2_lut_rep_399.init = 16'h6666;
    LUT4 i2_4_lut_then_4_lut (.A(ss[3]), .B(n21498), .C(ss[1]), .D(ss[0]), 
         .Z(n21505)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+!(C (D)))) */ ;
    defparam i2_4_lut_then_4_lut.init = 16'hefdf;
    LUT4 i2_4_lut_else_4_lut (.A(ss[3]), .B(n21498), .C(ss[1]), .D(ss[0]), 
         .Z(n21504)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i2_4_lut_else_4_lut.init = 16'hefd0;
    CCU2D add_15124_7 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18529), .COUT(n18530));
    defparam add_15124_7.INIT0 = 16'h0aaa;
    defparam add_15124_7.INIT1 = 16'hf555;
    defparam add_15124_7.INJECT1_0 = "NO";
    defparam add_15124_7.INJECT1_1 = "NO";
    CCU2D add_15134_21 (.A0(speed_set_m2[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18471), .S1(n42));
    defparam add_15134_21.INIT0 = 16'h5555;
    defparam add_15134_21.INIT1 = 16'h0000;
    defparam add_15134_21.INJECT1_0 = "NO";
    defparam add_15134_21.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(n1322[5]), .B(n1322[8]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 mux_1222_i10_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[9]), 
         .D(speed_set_m3[9]), .Z(n5365)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_then_4_lut (.A(n22216), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21508)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_else_4_lut (.A(n22216), .B(ss[1]), .C(ss[2]), .D(ss[3]), 
         .Z(n21507)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0100;
    CCU2D add_15124_5 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18528), .COUT(n18529));
    defparam add_15124_5.INIT0 = 16'h0aaa;
    defparam add_15124_5.INIT1 = 16'h0aaa;
    defparam add_15124_5.INJECT1_0 = "NO";
    defparam add_15124_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_392 (.A(ss[0]), .B(ss[2]), .Z(n21493)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_392.init = 16'h8888;
    LUT4 i1_2_lut_rep_361_3_lut (.A(ss[0]), .B(ss[2]), .C(ss[1]), .Z(n21462)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_361_3_lut.init = 16'h8080;
    LUT4 i11774_2_lut_3_lut_4_lut (.A(n22216), .B(n21458), .C(clk_N_875_enable_392), 
         .D(ss[1]), .Z(n14360)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11774_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i11802_2_lut_3_lut_4_lut (.A(n22216), .B(n21458), .C(clk_N_875_enable_303), 
         .D(ss[1]), .Z(n14388)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i11802_2_lut_3_lut_4_lut.init = 16'he0f0;
    FD1S3AX multOut_i0 (.D(multOut_28__N_1412[0]), .CK(clk_N_875), .Q(multOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i0.GSR = "ENABLED";
    CCU2D add_15124_3 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18527), .COUT(n18528));
    defparam add_15124_3.INIT0 = 16'hf555;
    defparam add_15124_3.INIT1 = 16'hf555;
    defparam add_15124_3.INJECT1_0 = "NO";
    defparam add_15124_3.INJECT1_1 = "NO";
    CCU2D add_15124_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[4]), .B1(speed_set_m2[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18527));
    defparam add_15124_1.INIT0 = 16'hF000;
    defparam add_15124_1.INIT1 = 16'ha666;
    defparam add_15124_1.INJECT1_0 = "NO";
    defparam add_15124_1.INJECT1_1 = "NO";
    CCU2D add_15125_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18526), 
          .S0(n1068));
    defparam add_15125_cout.INIT0 = 16'h0000;
    defparam add_15125_cout.INIT1 = 16'h0000;
    defparam add_15125_cout.INJECT1_0 = "NO";
    defparam add_15125_cout.INJECT1_1 = "NO";
    CCU2D add_15134_19 (.A0(speed_set_m2[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18470), .COUT(n18471));
    defparam add_15134_19.INIT0 = 16'hf555;
    defparam add_15134_19.INIT1 = 16'hf555;
    defparam add_15134_19.INJECT1_0 = "NO";
    defparam add_15134_19.INJECT1_1 = "NO";
    CCU2D add_15134_17 (.A0(speed_set_m2[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18469), .COUT(n18470));
    defparam add_15134_17.INIT0 = 16'hf555;
    defparam add_15134_17.INIT1 = 16'hf555;
    defparam add_15134_17.INJECT1_0 = "NO";
    defparam add_15134_17.INJECT1_1 = "NO";
    CCU2D add_15125_22 (.A0(addOut[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18525), .COUT(n18526));
    defparam add_15125_22.INIT0 = 16'h5555;
    defparam add_15125_22.INIT1 = 16'hf555;
    defparam add_15125_22.INJECT1_0 = "NO";
    defparam add_15125_22.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_11 (.A0(multOut[9]), .B0(n16420), .C0(addOut[9]), 
          .D0(addIn2_28__N_1441[9]), .A1(multOut[10]), .B1(n16420), .C1(addOut[10]), 
          .D1(addIn2_28__N_1441[10]), .CIN(n18411), .COUT(n18412), .S0(n121[9]), 
          .S1(n121[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_11.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_11.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_11.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_11.INJECT1_1 = "NO";
    CCU2D add_15134_15 (.A0(speed_set_m2[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18468), .COUT(n18469));
    defparam add_15134_15.INIT0 = 16'hf555;
    defparam add_15134_15.INIT1 = 16'hf555;
    defparam add_15134_15.INJECT1_0 = "NO";
    defparam add_15134_15.INJECT1_1 = "NO";
    CCU2D add_15125_20 (.A0(addOut[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18524), .COUT(n18525));
    defparam add_15125_20.INIT0 = 16'h5555;
    defparam add_15125_20.INIT1 = 16'h5555;
    defparam add_15125_20.INJECT1_0 = "NO";
    defparam add_15125_20.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n1322[3]), .B(n1322[2]), .C(n1322[1]), .D(n1322[0]), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'haaa8;
    LUT4 mux_1222_i6_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[5]), 
         .D(speed_set_m3[5]), .Z(n5357)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1222_i17_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[16]), 
         .D(speed_set_m3[16]), .Z(n5379)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i17_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_1206_3 (.A0(n1301[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1301[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18226), 
          .COUT(n18227), .S0(n2281[1]), .S1(n2281[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1206_3.INIT0 = 16'hf555;
    defparam add_1206_3.INIT1 = 16'hf555;
    defparam add_1206_3.INJECT1_0 = "NO";
    defparam add_1206_3.INJECT1_1 = "NO";
    CCU2D add_15134_13 (.A0(speed_set_m2[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18467), .COUT(n18468));
    defparam add_15134_13.INIT0 = 16'hf555;
    defparam add_15134_13.INIT1 = 16'hf555;
    defparam add_15134_13.INJECT1_0 = "NO";
    defparam add_15134_13.INJECT1_1 = "NO";
    CCU2D add_15125_18 (.A0(addOut[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18523), .COUT(n18524));
    defparam add_15125_18.INIT0 = 16'h5555;
    defparam add_15125_18.INIT1 = 16'h5555;
    defparam add_15125_18.INJECT1_0 = "NO";
    defparam add_15125_18.INJECT1_1 = "NO";
    LUT4 i9227_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[2]), .C(ss[3]), .D(ss[1]), 
         .Z(n15)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i9227_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_rep_393 (.A(n22216), .B(n22209), .Z(n21494)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_393.init = 16'hbbbb;
    LUT4 i1_3_lut (.A(n1322[15]), .B(n2293[8]), .C(n30), .Z(n19107)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[4] 360[11])
    defparam i1_3_lut.init = 16'h8a8a;
    CCU2D add_15125_16 (.A0(addOut[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18522), .COUT(n18523));
    defparam add_15125_16.INIT0 = 16'h5aaa;
    defparam add_15125_16.INIT1 = 16'h5555;
    defparam add_15125_16.INJECT1_0 = "NO";
    defparam add_15125_16.INJECT1_1 = "NO";
    CCU2D add_1206_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1301[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18226), 
          .S1(n2281[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1206_1.INIT0 = 16'hF000;
    defparam add_1206_1.INIT1 = 16'h0aaa;
    defparam add_1206_1.INJECT1_0 = "NO";
    defparam add_1206_1.INJECT1_1 = "NO";
    LUT4 mux_1222_i15_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[14]), 
         .D(speed_set_m3[14]), .Z(n5375)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_adj_42 (.A(n1322[15]), .B(n2293[7]), .C(n30), .Z(n19101)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[4] 360[11])
    defparam i1_3_lut_adj_42.init = 16'h8a8a;
    CCU2D addOut_2126_add_4_9 (.A0(multOut[7]), .B0(n16420), .C0(addOut[7]), 
          .D0(addIn2_28__N_1441[7]), .A1(multOut[8]), .B1(n16420), .C1(addOut[8]), 
          .D1(addIn2_28__N_1441[8]), .CIN(n18410), .COUT(n18411), .S0(n121[7]), 
          .S1(n121[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_9.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_9.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_9.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_9.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut (.A(n21407), .B(n21406), .C(n21410), .D(subIn1_24__N_1342), 
         .Z(n11585)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_189_i19_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[18]), 
         .Z(intgOut0_28__N_1629[18])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i19_3_lut_3_lut.init = 16'hbaba;
    CCU2D addOut_2126_add_4_7 (.A0(multOut[5]), .B0(n16420), .C0(addOut[5]), 
          .D0(addIn2_28__N_1441[5]), .A1(multOut[6]), .B1(n16420), .C1(addOut[6]), 
          .D1(addIn2_28__N_1441[6]), .CIN(n18409), .COUT(n18410), .S0(n121[5]), 
          .S1(n121[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_7.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_7.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_7.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_7.INJECT1_1 = "NO";
    FD1P3AX Out0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_97), .CK(clk_N_875), 
            .Q(Out0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i0.GSR = "ENABLED";
    FD1P3AX Out1_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i0.GSR = "ENABLED";
    FD1P3AX Out2_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i0.GSR = "ENABLED";
    FD1P3AX Out3_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i0.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i0.GSR = "DISABLED";
    FD1S3IX ss_i2 (.D(n14), .CK(clk_N_875), .CD(ss[4]), .Q(ss[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i2.GSR = "ENABLED";
    FD1P3AX backOut3_i0_i0 (.D(Out3_28__N_1174[0]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i0.GSR = "DISABLED";
    FD1S3AX subOut_i0 (.D(\subOut_24__N_1369[0] ), .CK(clk_N_875), .Q(subOut[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i0.GSR = "ENABLED";
    CCU2D add_15125_14 (.A0(addOut[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18521), .COUT(n18522));
    defparam add_15125_14.INIT0 = 16'h5aaa;
    defparam add_15125_14.INIT1 = 16'h5555;
    defparam add_15125_14.INJECT1_0 = "NO";
    defparam add_15125_14.INJECT1_1 = "NO";
    LUT4 mux_1222_i2_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[1]), 
         .D(speed_set_m3[1]), .Z(n5349)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1222_i11_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[10]), 
         .D(speed_set_m3[10]), .Z(n5367)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i11_3_lut_4_lut.init = 16'hfb40;
    CCU2D addOut_2126_add_4_5 (.A0(multOut[3]), .B0(n16420), .C0(addOut[3]), 
          .D0(addIn2_28__N_1441[3]), .A1(multOut[4]), .B1(n16420), .C1(addOut[4]), 
          .D1(addIn2_28__N_1441[4]), .CIN(n18408), .COUT(n18409), .S0(n121[3]), 
          .S1(n121[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_5.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_5.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_5.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_5.INJECT1_1 = "NO";
    CCU2D add_15134_11 (.A0(speed_set_m2[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18466), .COUT(n18467));
    defparam add_15134_11.INIT0 = 16'hf555;
    defparam add_15134_11.INIT1 = 16'hf555;
    defparam add_15134_11.INJECT1_0 = "NO";
    defparam add_15134_11.INJECT1_1 = "NO";
    CCU2D add_15125_12 (.A0(addOut[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18520), .COUT(n18521));
    defparam add_15125_12.INIT0 = 16'h5555;
    defparam add_15125_12.INIT1 = 16'h5aaa;
    defparam add_15125_12.INJECT1_0 = "NO";
    defparam add_15125_12.INJECT1_1 = "NO";
    CCU2D add_15134_9 (.A0(speed_set_m2[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18465), .COUT(n18466));
    defparam add_15134_9.INIT0 = 16'hf555;
    defparam add_15134_9.INIT1 = 16'hf555;
    defparam add_15134_9.INJECT1_0 = "NO";
    defparam add_15134_9.INJECT1_1 = "NO";
    LUT4 mux_1222_i7_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[6]), 
         .D(speed_set_m3[6]), .Z(n5359)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1222_i3_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[2]), 
         .D(speed_set_m3[2]), .Z(n5351)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13900_2_lut_rep_309 (.A(n16496), .B(n42), .Z(n21410)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13900_2_lut_rep_309.init = 16'heeee;
    LUT4 i1_4_lut_4_lut (.A(n22216), .B(n21463), .C(n21462), .D(ss[3]), 
         .Z(clk_N_875_enable_181)) /* synthesis lut_function=(A (B)+!A (C (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_4_lut_4_lut.init = 16'hd888;
    CCU2D add_15134_7 (.A0(speed_set_m2[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18464), .COUT(n18465));
    defparam add_15134_7.INIT0 = 16'hf555;
    defparam add_15134_7.INIT1 = 16'hf555;
    defparam add_15134_7.INJECT1_0 = "NO";
    defparam add_15134_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_363_3_lut (.A(n22216), .B(ss[2]), .C(ss[3]), .Z(n21464)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_363_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_366_3_lut (.A(n22216), .B(n22209), .C(ss[3]), .Z(n21467)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_366_3_lut.init = 16'hfbfb;
    CCU2D add_15125_10 (.A0(addOut[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18519), .COUT(n18520));
    defparam add_15125_10.INIT0 = 16'h5aaa;
    defparam add_15125_10.INIT1 = 16'h5aaa;
    defparam add_15125_10.INJECT1_0 = "NO";
    defparam add_15125_10.INJECT1_1 = "NO";
    LUT4 equal_112_i9_2_lut_3_lut_4_lut (.A(n22216), .B(n22209), .C(n6), 
         .D(ss[3]), .Z(n9)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam equal_112_i9_2_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 equal_133_i9_2_lut_3_lut_4_lut (.A(n22216), .B(ss[2]), .C(n21495), 
         .D(ss[3]), .Z(n9_adj_2327)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam equal_133_i9_2_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 ss_4__I_0_351_i6_2_lut_rep_394 (.A(ss[0]), .B(ss[1]), .Z(n21495)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(164[29:36])
    defparam ss_4__I_0_351_i6_2_lut_rep_394.init = 16'hbbbb;
    CCU2D addOut_2126_add_4_3 (.A0(multOut[1]), .B0(n16420), .C0(addOut[1]), 
          .D0(addIn2_28__N_1441[1]), .A1(multOut[2]), .B1(n16420), .C1(addOut[2]), 
          .D1(addIn2_28__N_1441[2]), .CIN(n18407), .COUT(n18408), .S0(n121[1]), 
          .S1(n121[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_3.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_3.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_3.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_43 (.A(n1322[15]), .B(n2293[6]), .C(n30), .Z(n1458[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_43.init = 16'h8a8a;
    LUT4 i17204_2_lut_rep_302_3_lut_3_lut_4_lut (.A(n16496), .B(n42), .C(subIn1_24__N_1342), 
         .D(n35), .Z(n21403)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)))) */ ;
    defparam i17204_2_lut_rep_302_3_lut_3_lut_4_lut.init = 16'h11f1;
    LUT4 i1_4_lut_4_lut_adj_44 (.A(n22216), .B(n21463), .C(n19679), .D(ss[1]), 
         .Z(clk_N_875_enable_97)) /* synthesis lut_function=(A (B)+!A !(C+(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_4_lut_4_lut_adj_44.init = 16'h888d;
    CCU2D add_15125_8 (.A0(addOut[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18518), .COUT(n18519));
    defparam add_15125_8.INIT0 = 16'h5555;
    defparam add_15125_8.INIT1 = 16'h5aaa;
    defparam add_15125_8.INJECT1_0 = "NO";
    defparam add_15125_8.INJECT1_1 = "NO";
    LUT4 mux_189_i17_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[16]), 
         .Z(intgOut0_28__N_1629[16])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i17_3_lut_3_lut.init = 16'hbaba;
    CCU2D add_1209_11 (.A0(n1364[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18338), 
          .S0(n2317[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1209_11.INIT0 = 16'hf555;
    defparam add_1209_11.INIT1 = 16'h0000;
    defparam add_1209_11.INJECT1_0 = "NO";
    defparam add_1209_11.INJECT1_1 = "NO";
    CCU2D add_1209_9 (.A0(n1364[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1364[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18337), 
          .COUT(n18338), .S0(n2317[7]), .S1(n2317[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1209_9.INIT0 = 16'hf555;
    defparam add_1209_9.INIT1 = 16'hf555;
    defparam add_1209_9.INJECT1_0 = "NO";
    defparam add_1209_9.INJECT1_1 = "NO";
    CCU2D add_1212_7 (.A0(n5443), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5445), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18233), 
          .COUT(n18234), .S0(n2373[5]), .S1(n2373[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_7.INIT0 = 16'hf555;
    defparam add_1212_7.INIT1 = 16'hf555;
    defparam add_1212_7.INJECT1_0 = "NO";
    defparam add_1212_7.INJECT1_1 = "NO";
    CCU2D add_15125_6 (.A0(addOut[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18517), .COUT(n18518));
    defparam add_15125_6.INIT0 = 16'h5555;
    defparam add_15125_6.INIT1 = 16'h5555;
    defparam add_15125_6.INJECT1_0 = "NO";
    defparam add_15125_6.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_45 (.A(n1322[15]), .B(n2293[5]), .C(n30), .Z(n1458[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_45.init = 16'h8a8a;
    LUT4 mux_1221_i14_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m4[13]), .Z(n5415)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_4_lut_adj_46 (.A(n22216), .B(n21463), .C(n19679), .D(ss[1]), 
         .Z(clk_N_875_enable_153)) /* synthesis lut_function=(A (B)+!A !(C+!(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_4_lut_4_lut_adj_46.init = 16'h8d88;
    LUT4 i1_4_lut_4_lut_adj_47 (.A(n22216), .B(n21463), .C(n21474), .D(n11644), 
         .Z(clk_N_875_enable_125)) /* synthesis lut_function=(A (B)+!A (C (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_4_lut_4_lut_adj_47.init = 16'hd888;
    LUT4 i1_2_lut_rep_397 (.A(n22216), .B(n22209), .Z(n21498)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_397.init = 16'heeee;
    FD1S3IX ss_i3 (.D(n15), .CK(clk_N_875), .CD(ss[4]), .Q(ss[3]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i3.GSR = "ENABLED";
    FD1P3IX intgOut3_i0 (.D(addOut[0]), .SP(clk_N_875_enable_303), .CD(n14382), 
            .CK(clk_N_875), .Q(intgOut3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i0.GSR = "ENABLED";
    LUT4 i11815_4_lut (.A(clk_N_875_enable_391), .B(n21463), .C(n30), 
         .D(n1322[15]), .Z(n14419)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11815_4_lut.init = 16'h8aaa;
    LUT4 i1_3_lut_adj_48 (.A(n1322[15]), .B(n2293[3]), .C(n30), .Z(n1458[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_48.init = 16'h8a8a;
    LUT4 mux_136_i6_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[5]), 
         .D(backOut1[5]), .Z(n588[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i22_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[21]), 
         .D(backOut1[21]), .Z(n588[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1221_i8_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m4[7]), .Z(n5403)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i4_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[3]), 
         .D(backOut1[3]), .Z(n588[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_365_3_lut (.A(n22216), .B(ss[2]), .C(ss[3]), .Z(n21466)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_365_3_lut.init = 16'hfefe;
    LUT4 i13934_2_lut_3_lut_4_lut (.A(n16496), .B(n42), .C(n49), .D(n15773), 
         .Z(n16542)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i13934_2_lut_3_lut_4_lut.init = 16'heee0;
    LUT4 mux_189_i16_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[15]), 
         .Z(intgOut0_28__N_1629[15])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i16_3_lut_3_lut.init = 16'hbaba;
    LUT4 i1_2_lut_rep_370_3_lut (.A(n22216), .B(n22209), .C(ss[3]), .Z(n21471)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam i1_2_lut_rep_370_3_lut.init = 16'hefef;
    LUT4 mux_136_i3_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[2]), 
         .D(backOut1[2]), .Z(n588[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i1_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[0]), 
         .D(backOut1[0]), .Z(n588[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_189_i15_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[14]), 
         .Z(intgOut0_28__N_1629[14])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i15_3_lut_3_lut.init = 16'hbaba;
    LUT4 i13126_2_lut_rep_398 (.A(n22216), .B(ss[3]), .Z(n21499)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13126_2_lut_rep_398.init = 16'heeee;
    LUT4 i1_2_lut_rep_369_3_lut_4_lut (.A(n22216), .B(ss[3]), .C(ss[1]), 
         .D(ss[0]), .Z(n21470)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_rep_369_3_lut_4_lut.init = 16'h0110;
    LUT4 mux_136_i29_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[28]), 
         .D(backOut1[28]), .Z(n588[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i29_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15137_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18225), 
          .S0(n35));
    defparam add_15137_cout.INIT0 = 16'h0000;
    defparam add_15137_cout.INIT1 = 16'h0000;
    defparam add_15137_cout.INJECT1_0 = "NO";
    defparam add_15137_cout.INJECT1_1 = "NO";
    CCU2D add_15134_5 (.A0(speed_set_m2[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18463), .COUT(n18464));
    defparam add_15134_5.INIT0 = 16'hf555;
    defparam add_15134_5.INIT1 = 16'hf555;
    defparam add_15134_5.INJECT1_0 = "NO";
    defparam add_15134_5.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(multOut[0]), .B1(n16420), .C1(addOut[0]), 
          .D1(addIn2_28__N_1441[0]), .COUT(n18407), .S1(n121[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_1.INIT0 = 16'hF000;
    defparam addOut_2126_add_4_1.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_1.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_1.INJECT1_1 = "NO";
    CCU2D add_15137_21 (.A0(speed_set_m1[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18224), .COUT(n18225));
    defparam add_15137_21.INIT0 = 16'hf555;
    defparam add_15137_21.INIT1 = 16'h5555;
    defparam add_15137_21.INJECT1_0 = "NO";
    defparam add_15137_21.INJECT1_1 = "NO";
    LUT4 mux_136_i23_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[22]), 
         .D(backOut1[22]), .Z(n588[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i5_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[4]), 
         .D(backOut1[4]), .Z(n588[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i28_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[27]), 
         .D(backOut1[27]), .Z(n588[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i27_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[26]), 
         .D(backOut1[26]), .Z(n588[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i27_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15125_4 (.A0(addOut[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18516), .COUT(n18517));
    defparam add_15125_4.INIT0 = 16'h5aaa;
    defparam add_15125_4.INIT1 = 16'h5aaa;
    defparam add_15125_4.INJECT1_0 = "NO";
    defparam add_15125_4.INJECT1_1 = "NO";
    CCU2D add_15134_3 (.A0(speed_set_m2[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18462), .COUT(n18463));
    defparam add_15134_3.INIT0 = 16'hf555;
    defparam add_15134_3.INIT1 = 16'hf555;
    defparam add_15134_3.INJECT1_0 = "NO";
    defparam add_15134_3.INJECT1_1 = "NO";
    CCU2D add_15134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m2[0]), .B1(speed_set_m2[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18462));
    defparam add_15134_1.INIT0 = 16'hF000;
    defparam add_15134_1.INIT1 = 16'ha666;
    defparam add_15134_1.INJECT1_0 = "NO";
    defparam add_15134_1.INJECT1_1 = "NO";
    LUT4 mux_136_i26_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[25]), 
         .D(backOut1[25]), .Z(n588[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i25_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[24]), 
         .D(backOut1[24]), .Z(n588[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i24_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[23]), 
         .D(backOut1[23]), .Z(n588[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_189_i11_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[10]), 
         .Z(intgOut0_28__N_1629[10])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i11_3_lut_3_lut.init = 16'hbaba;
    LUT4 mux_136_i2_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[1]), 
         .D(backOut1[1]), .Z(n588[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_189_i10_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[9]), 
         .Z(intgOut0_28__N_1629[9])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i10_3_lut_3_lut.init = 16'hbaba;
    LUT4 mux_136_i7_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[6]), 
         .D(backOut1[6]), .Z(n588[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i8_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[7]), 
         .D(backOut1[7]), .Z(n588[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i9_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[8]), 
         .D(backOut1[8]), .Z(n588[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i10_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[9]), 
         .D(backOut1[9]), .Z(n588[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i11_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[10]), 
         .D(backOut1[10]), .Z(n588[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_1221_i13_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m4[12]), .Z(n5413)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_136_i12_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[11]), 
         .D(backOut1[11]), .Z(n588[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i13_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[12]), 
         .D(backOut1[12]), .Z(n588[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i14_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[13]), 
         .D(backOut1[13]), .Z(n588[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i15_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[14]), 
         .D(backOut1[14]), .Z(n588[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i16_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[15]), 
         .D(backOut1[15]), .Z(n588[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i17_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[16]), 
         .D(backOut1[16]), .Z(n588[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i18_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[17]), 
         .D(backOut1[17]), .Z(n588[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i19_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[18]), 
         .D(backOut1[18]), .Z(n588[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_136_i20_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[19]), 
         .D(backOut1[19]), .Z(n588[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_adj_49 (.A(n1301[15]), .B(n2281[9]), .C(n9_adj_2328), 
         .Z(n1414[9])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_49.init = 16'h8a8a;
    CCU2D add_15137_19 (.A0(speed_set_m1[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18223), .COUT(n18224));
    defparam add_15137_19.INIT0 = 16'hf555;
    defparam add_15137_19.INIT1 = 16'hf555;
    defparam add_15137_19.INJECT1_0 = "NO";
    defparam add_15137_19.INJECT1_1 = "NO";
    CCU2D add_15137_17 (.A0(speed_set_m1[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18222), .COUT(n18223));
    defparam add_15137_17.INIT0 = 16'hf555;
    defparam add_15137_17.INIT1 = 16'hf555;
    defparam add_15137_17.INJECT1_0 = "NO";
    defparam add_15137_17.INJECT1_1 = "NO";
    LUT4 mux_136_i21_3_lut_4_lut (.A(n21473), .B(n21471), .C(backOut0[20]), 
         .D(backOut1[20]), .Z(n588[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(173[9:17])
    defparam mux_136_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5_4_lut (.A(n9_adj_2329), .B(n1301[10]), .C(n8_adj_2330), .D(n1301[11]), 
         .Z(n9_adj_2328)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i3_2_lut (.A(n1301[14]), .B(n1301[13]), .Z(n9_adj_2329)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    CCU2D add_15127_29 (.A0(addOut[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18461), 
          .S1(n3840));
    defparam add_15127_29.INIT0 = 16'h5aaa;
    defparam add_15127_29.INIT1 = 16'h0000;
    defparam add_15127_29.INJECT1_0 = "NO";
    defparam add_15127_29.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n1301[9]), .B(n1301[12]), .C(n10_adj_2331), .D(n1301[7]), 
         .Z(n8_adj_2330)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'hccc8;
    CCU2D add_15137_15 (.A0(speed_set_m1[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18221), .COUT(n18222));
    defparam add_15137_15.INIT0 = 16'hf555;
    defparam add_15137_15.INIT1 = 16'hf555;
    defparam add_15137_15.INJECT1_0 = "NO";
    defparam add_15137_15.INJECT1_1 = "NO";
    LUT4 i4_4_lut_adj_50 (.A(n1301[6]), .B(n8_adj_2332), .C(n1301[4]), 
         .D(n4_adj_2333), .Z(n10_adj_2331)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_50.init = 16'hfeee;
    CCU2D add_15137_13 (.A0(speed_set_m1[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18220), .COUT(n18221));
    defparam add_15137_13.INIT0 = 16'hf555;
    defparam add_15137_13.INIT1 = 16'hf555;
    defparam add_15137_13.INJECT1_0 = "NO";
    defparam add_15137_13.INJECT1_1 = "NO";
    LUT4 i2_2_lut_adj_51 (.A(n1301[5]), .B(n1301[8]), .Z(n8_adj_2332)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_51.init = 16'heeee;
    LUT4 i1_4_lut_adj_52 (.A(n1301[3]), .B(n1301[2]), .C(n1301[1]), .D(n1301[0]), 
         .Z(n4_adj_2333)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_52.init = 16'haaa8;
    CCU2D add_15137_3 (.A0(speed_set_m1[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18215), .COUT(n18216));
    defparam add_15137_3.INIT0 = 16'hf555;
    defparam add_15137_3.INIT1 = 16'hf555;
    defparam add_15137_3.INJECT1_0 = "NO";
    defparam add_15137_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_53 (.A(n1301[15]), .B(n2281[8]), .C(n9_adj_2328), 
         .Z(n1414[8])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_53.init = 16'h8a8a;
    LUT4 mux_139_i2_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[1]), 
         .D(n648[1]), .Z(n678[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i2_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15137_7 (.A0(speed_set_m1[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18217), .COUT(n18218));
    defparam add_15137_7.INIT0 = 16'hf555;
    defparam add_15137_7.INIT1 = 16'hf555;
    defparam add_15137_7.INJECT1_0 = "NO";
    defparam add_15137_7.INJECT1_1 = "NO";
    LUT4 mux_139_i3_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[2]), 
         .D(n648[2]), .Z(n678[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i3_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15137_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18215));
    defparam add_15137_1.INIT0 = 16'hF000;
    defparam add_15137_1.INIT1 = 16'h0aaa;
    defparam add_15137_1.INJECT1_0 = "NO";
    defparam add_15137_1.INJECT1_1 = "NO";
    FD1S3AY ss_i4 (.D(n19674), .CK(clk_N_875), .Q(ss[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i4.GSR = "ENABLED";
    LUT4 i1_3_lut_adj_54 (.A(n1301[15]), .B(n2281[7]), .C(n9_adj_2328), 
         .Z(n1414[7])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_54.init = 16'h8a8a;
    CCU2D add_15137_11 (.A0(speed_set_m1[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18219), .COUT(n18220));
    defparam add_15137_11.INIT0 = 16'hf555;
    defparam add_15137_11.INIT1 = 16'hf555;
    defparam add_15137_11.INJECT1_0 = "NO";
    defparam add_15137_11.INJECT1_1 = "NO";
    CCU2D add_15137_5 (.A0(speed_set_m1[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18216), .COUT(n18217));
    defparam add_15137_5.INIT0 = 16'hf555;
    defparam add_15137_5.INIT1 = 16'hf555;
    defparam add_15137_5.INJECT1_0 = "NO";
    defparam add_15137_5.INJECT1_1 = "NO";
    LUT4 mux_139_i19_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[18]), 
         .D(n648[18]), .Z(n678[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i19_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15137_9 (.A0(speed_set_m1[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18218), .COUT(n18219));
    defparam add_15137_9.INIT0 = 16'hf555;
    defparam add_15137_9.INIT1 = 16'hf555;
    defparam add_15137_9.INJECT1_0 = "NO";
    defparam add_15137_9.INJECT1_1 = "NO";
    CCU2D add_15125_2 (.A0(addOut[7]), .B0(addOut[6]), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18516));
    defparam add_15125_2.INIT0 = 16'h7000;
    defparam add_15125_2.INIT1 = 16'h5555;
    defparam add_15125_2.INJECT1_0 = "NO";
    defparam add_15125_2.INJECT1_1 = "NO";
    LUT4 mux_139_i18_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[17]), 
         .D(n648[17]), .Z(n678[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i13_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[12]), 
         .D(n648[12]), .Z(n678[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_adj_55 (.A(n1301[15]), .B(n2281[6]), .C(n9_adj_2328), 
         .Z(n1414[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_55.init = 16'h8a8a;
    LUT4 i1_3_lut_adj_56 (.A(n1301[15]), .B(n2281[5]), .C(n9_adj_2328), 
         .Z(n1414[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_56.init = 16'h8a8a;
    LUT4 i3382_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m2[9]), .Z(n5884)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3382_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i11_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[10]), 
         .D(n648[10]), .Z(n678[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11806_4_lut (.A(clk_N_875_enable_391), .B(n1301[15]), .C(n9_adj_2328), 
         .D(n21463), .Z(n14410)) /* synthesis lut_function=(A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11806_4_lut.init = 16'haa2a;
    LUT4 mux_139_i10_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[9]), 
         .D(n648[9]), .Z(n678[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_adj_57 (.A(n1301[15]), .B(n2281[3]), .C(n9_adj_2328), 
         .Z(n1414[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_57.init = 16'h8a8a;
    LUT4 mux_139_i4_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[3]), 
         .D(n648[3]), .Z(n678[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_189_i8_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[7]), 
         .Z(intgOut0_28__N_1629[7])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i8_3_lut_3_lut.init = 16'hbaba;
    FD1P3AX dirout_m2_347 (.D(subIn1_24__N_1534), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m2));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m2_347.GSR = "DISABLED";
    FD1P3AX dirout_m3_348 (.D(dirout_m3_N_1949), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m3));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m3_348.GSR = "DISABLED";
    FD1P3AX dirout_m1_346 (.D(subIn1_24__N_1347), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m1));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m1_346.GSR = "DISABLED";
    FD1P3AX dirout_m4_349 (.D(dirout_m4_N_1952), .SP(clk_N_875_enable_391), 
            .CK(clk_N_875), .Q(dir_m4));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dirout_m4_349.GSR = "DISABLED";
    LUT4 mux_139_i25_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[24]), 
         .D(n648[24]), .Z(n678[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i25_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX backOut1_i0_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i28.GSR = "DISABLED";
    LUT4 mux_139_i24_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[23]), 
         .D(n648[23]), .Z(n678[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i20_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[19]), 
         .D(n648[19]), .Z(n678[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i20_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_15127_27 (.A0(addOut[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18460), .COUT(n18461));
    defparam add_15127_27.INIT0 = 16'h0aaa;
    defparam add_15127_27.INIT1 = 16'h0aaa;
    defparam add_15127_27.INJECT1_0 = "NO";
    defparam add_15127_27.INJECT1_1 = "NO";
    FD1P3AX backOut1_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i25.GSR = "DISABLED";
    CCU2D add_223_17 (.A0(Out3[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18273), 
          .S0(n1364[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_17.INIT0 = 16'h5aaa;
    defparam add_223_17.INIT1 = 16'h0000;
    defparam add_223_17.INJECT1_0 = "NO";
    defparam add_223_17.INJECT1_1 = "NO";
    FD1P3AX backOut1_i0_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i6.GSR = "DISABLED";
    LUT4 mux_139_i29_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[28]), 
         .D(n648[28]), .Z(n678[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i29_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX backOut1_i0_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut1_i0_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_41), 
            .CK(clk_N_875), .Q(backOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut1_i0_i1.GSR = "DISABLED";
    LUT4 mux_139_i8_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[7]), 
         .D(n648[7]), .Z(n678[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i17_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[16]), 
         .D(n648[16]), .Z(n678[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i14_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[13]), 
         .D(n648[13]), .Z(n678[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i12_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[11]), 
         .D(n648[11]), .Z(n678[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i9_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[8]), 
         .D(n648[8]), .Z(n678[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i5_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[4]), 
         .D(n648[4]), .Z(n678[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3145_3_lut (.A(n3840), .B(n1068), .C(addOut[28]), .Z(intgOut0_28__N_1629[28])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3145_3_lut.init = 16'h3232;
    LUT4 mux_139_i15_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[14]), 
         .D(n648[14]), .Z(n678[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i26_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[25]), 
         .D(n648[25]), .Z(n678[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i23_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[22]), 
         .D(n648[22]), .Z(n678[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i16_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[15]), 
         .D(n648[15]), .Z(n678[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3054_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m2[0]), .Z(n5556)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3054_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i22_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[21]), 
         .D(n648[21]), .Z(n678[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i13_3_lut (.A(\speed_avg_m3[12] ), .B(\speed_avg_m2[12] ), 
         .C(n22204), .Z(subIn2_24__N_1535[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i13_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_58 (.A(n16258), .B(n19662), .C(n22216), .D(n21493), 
         .Z(clk_N_875_enable_69)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_58.init = 16'hc4c0;
    LUT4 mux_139_i27_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[26]), 
         .D(n648[26]), .Z(n678[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i6_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[5]), 
         .D(n648[5]), .Z(n678[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i7_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[6]), 
         .D(n648[6]), .Z(n678[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i28_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[27]), 
         .D(n648[27]), .Z(n678[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i21_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[20]), 
         .D(n648[20]), .Z(n678[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_139_i1_3_lut_4_lut (.A(n21473), .B(n21466), .C(intgOut0[0]), 
         .D(n648[0]), .Z(n678[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam mux_139_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13249_2_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[6]), .Z(intgOut0_28__N_1629[6])) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i13249_2_lut_3_lut.init = 16'hfefe;
    LUT4 i11779_3_lut_4_lut (.A(n1068), .B(n3840), .C(n21424), .D(clk_N_875_enable_303), 
         .Z(n14382)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i11779_3_lut_4_lut.init = 16'hfe00;
    LUT4 i3366_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m2[1]), .Z(n5868)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3366_3_lut_4_lut.init = 16'hfd20;
    LUT4 subIn2_24__I_25_i13_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[12] ), 
         .D(subIn2_24__N_1535[12]), .Z(subIn2_24__N_1348[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i10_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[9] ), 
         .D(subIn2_24__N_1535[9]), .Z(subIn2_24__N_1348[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i9_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[8] ), 
         .D(subIn2_24__N_1535[8]), .Z(subIn2_24__N_1348[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i9_3_lut_4_lut.init = 16'hfb40;
    FD1S3AX addOut_2126__i0 (.D(n121[0]), .CK(clk_N_875), .Q(addOut[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i0.GSR = "ENABLED";
    AND2 AND2_t64 (.A(subOut[0]), .B(multIn2[0]), .Z(multOut_28__N_1412[0])) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1256[10:66])
    AND2 AND2_t61 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1262[10:66])
    AND2 AND2_t58 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1268[10:66])
    AND2 AND2_t55 (.A(subOut[0]), .B(multIn2[3]), .Z(mult_29s_25s_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1274[10:66])
    AND2 AND2_t52 (.A(subOut[0]), .B(multIn2[9]), .Z(mult_29s_25s_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1280[10:66])
    AND2 AND2_t49 (.A(subOut[0]), .B(multIn2[11]), .Z(mult_29s_25s_0_pp_5_10)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1286[10:68])
    AND2 AND2_t46 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_6_12)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1292[10:68])
    AND2 AND2_t43 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_7_14)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1298[10:68])
    AND2 AND2_t40 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_8_16)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1304[10:68])
    AND2 AND2_t37 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_9_18)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1310[10:68])
    AND2 AND2_t34 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_10_20)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1316[10:69])
    AND2 AND2_t31 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_11_22)) /* synthesis syn_instantiated=1 */ ;   // mult_29s_25s.v(1322[10:69])
    ND2 ND2_t28 (.A(subOut[0]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t27 (.A(subOut[1]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_25)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t26 (.A(subOut[2]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t25 (.A(subOut[3]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_27)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    ND2 ND2_t24 (.A(subOut[4]), .B(GND_net), .Z(mult_29s_25s_0_pp_12_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i8_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[7] ), 
         .D(subIn2_24__N_1535[7]), .Z(subIn2_24__N_1348[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i4_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[3] ), 
         .D(subIn2_24__N_1535[3]), .Z(subIn2_24__N_1348[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i4_3_lut_4_lut.init = 16'hfb40;
    FADD2B mult_29s_25s_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_12 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_14 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_16 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_18 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_20 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_22 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_0_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_0_2), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_1_2), .CI(GND_net), .COUT(co_mult_29s_25s_0_0_1), 
           .S1(multOut_28__N_1412[2])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_2 (.A0(mult_29s_25s_0_pp_0_3), .A1(mult_29s_25s_0_pp_0_4), 
           .B0(mult_29s_25s_0_pp_1_3), .B1(mult_29s_25s_0_pp_1_4), .CI(co_mult_29s_25s_0_0_1), 
           .COUT(co_mult_29s_25s_0_0_2), .S0(multOut_28__N_1412[3]), .S1(s_mult_29s_25s_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_3 (.A0(mult_29s_25s_0_pp_0_5), .A1(mult_29s_25s_0_pp_0_6), 
           .B0(mult_29s_25s_0_pp_1_5), .B1(mult_29s_25s_0_pp_1_6), .CI(co_mult_29s_25s_0_0_2), 
           .COUT(co_mult_29s_25s_0_0_3), .S0(s_mult_29s_25s_0_0_5), .S1(s_mult_29s_25s_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_4 (.A0(mult_29s_25s_0_pp_0_7), .A1(mult_29s_25s_0_pp_0_8), 
           .B0(mult_29s_25s_0_pp_1_7), .B1(mult_29s_25s_0_pp_1_8), .CI(co_mult_29s_25s_0_0_3), 
           .COUT(co_mult_29s_25s_0_0_4), .S0(s_mult_29s_25s_0_0_7), .S1(s_mult_29s_25s_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_5 (.A0(mult_29s_25s_0_pp_0_9), .A1(mult_29s_25s_0_pp_0_10), 
           .B0(mult_29s_25s_0_pp_1_9), .B1(mult_29s_25s_0_pp_1_10), .CI(co_mult_29s_25s_0_0_4), 
           .COUT(co_mult_29s_25s_0_0_5), .S0(s_mult_29s_25s_0_0_9), .S1(s_mult_29s_25s_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_6 (.A0(mult_29s_25s_0_pp_0_11), .A1(mult_29s_25s_0_pp_0_12), 
           .B0(mult_29s_25s_0_pp_1_11), .B1(mult_29s_25s_0_pp_1_12), .CI(co_mult_29s_25s_0_0_5), 
           .COUT(co_mult_29s_25s_0_0_6), .S0(s_mult_29s_25s_0_0_11), .S1(s_mult_29s_25s_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_7 (.A0(mult_29s_25s_0_pp_0_13), .A1(mult_29s_25s_0_pp_0_14), 
           .B0(mult_29s_25s_0_pp_1_13), .B1(mult_29s_25s_0_pp_1_14), .CI(co_mult_29s_25s_0_0_6), 
           .COUT(co_mult_29s_25s_0_0_7), .S0(s_mult_29s_25s_0_0_13), .S1(s_mult_29s_25s_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_8 (.A0(mult_29s_25s_0_pp_0_15), .A1(mult_29s_25s_0_pp_0_16), 
           .B0(mult_29s_25s_0_pp_1_15), .B1(mult_29s_25s_0_pp_1_16), .CI(co_mult_29s_25s_0_0_7), 
           .COUT(co_mult_29s_25s_0_0_8), .S0(s_mult_29s_25s_0_0_15), .S1(s_mult_29s_25s_0_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_9 (.A0(mult_29s_25s_0_pp_0_17), .A1(mult_29s_25s_0_pp_0_18), 
           .B0(mult_29s_25s_0_pp_1_17), .B1(mult_29s_25s_0_pp_1_18), .CI(co_mult_29s_25s_0_0_8), 
           .COUT(co_mult_29s_25s_0_0_9), .S0(s_mult_29s_25s_0_0_17), .S1(s_mult_29s_25s_0_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_10 (.A0(mult_29s_25s_0_pp_0_19), .A1(mult_29s_25s_0_pp_0_20), 
           .B0(mult_29s_25s_0_pp_1_19), .B1(mult_29s_25s_0_pp_1_20), .CI(co_mult_29s_25s_0_0_9), 
           .COUT(co_mult_29s_25s_0_0_10), .S0(s_mult_29s_25s_0_0_19), .S1(s_mult_29s_25s_0_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_11 (.A0(mult_29s_25s_0_pp_0_21), .A1(mult_29s_25s_0_pp_0_22), 
           .B0(mult_29s_25s_0_pp_1_21), .B1(mult_29s_25s_0_pp_1_22), .CI(co_mult_29s_25s_0_0_10), 
           .COUT(co_mult_29s_25s_0_0_11), .S0(s_mult_29s_25s_0_0_21), .S1(s_mult_29s_25s_0_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_12 (.A0(mult_29s_25s_0_pp_0_23), .A1(mult_29s_25s_0_pp_0_24), 
           .B0(mult_29s_25s_0_pp_1_23), .B1(mult_29s_25s_0_pp_1_24), .CI(co_mult_29s_25s_0_0_11), 
           .COUT(co_mult_29s_25s_0_0_12), .S0(s_mult_29s_25s_0_0_23), .S1(s_mult_29s_25s_0_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_13 (.A0(mult_29s_25s_0_pp_0_25), .A1(mult_29s_25s_0_pp_0_26), 
           .B0(mult_29s_25s_0_pp_1_25), .B1(mult_29s_25s_0_pp_1_26), .CI(co_mult_29s_25s_0_0_12), 
           .COUT(co_mult_29s_25s_0_0_13), .S0(s_mult_29s_25s_0_0_25), .S1(s_mult_29s_25s_0_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_0_14 (.A0(mult_29s_25s_0_pp_0_27), .A1(mult_29s_25s_0_pp_0_28), 
           .B0(mult_29s_25s_0_pp_1_27), .B1(mult_29s_25s_0_pp_1_28), .CI(co_mult_29s_25s_0_0_13), 
           .S0(s_mult_29s_25s_0_0_27), .S1(s_mult_29s_25s_0_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i20_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[19] ), 
         .D(\speed_avg_m2[19] ), .Z(subIn2_24__N_1348[19])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i20_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_mult_29s_25s_0_1_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_2_6), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_3_6), .CI(GND_net), .COUT(co_mult_29s_25s_0_1_1), 
           .S1(s_mult_29s_25s_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_2 (.A0(mult_29s_25s_0_pp_2_7), .A1(mult_29s_25s_0_pp_2_8), 
           .B0(mult_29s_25s_0_pp_3_7), .B1(mult_29s_25s_0_pp_3_8), .CI(co_mult_29s_25s_0_1_1), 
           .COUT(co_mult_29s_25s_0_1_2), .S0(s_mult_29s_25s_0_1_7), .S1(s_mult_29s_25s_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_3 (.A0(mult_29s_25s_0_pp_2_9), .A1(mult_29s_25s_0_pp_2_10), 
           .B0(mult_29s_25s_0_pp_3_9), .B1(mult_29s_25s_0_pp_3_10), .CI(co_mult_29s_25s_0_1_2), 
           .COUT(co_mult_29s_25s_0_1_3), .S0(s_mult_29s_25s_0_1_9), .S1(s_mult_29s_25s_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_4 (.A0(mult_29s_25s_0_pp_2_11), .A1(mult_29s_25s_0_pp_2_12), 
           .B0(mult_29s_25s_0_pp_3_11), .B1(mult_29s_25s_0_pp_3_12), .CI(co_mult_29s_25s_0_1_3), 
           .COUT(co_mult_29s_25s_0_1_4), .S0(s_mult_29s_25s_0_1_11), .S1(s_mult_29s_25s_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_5 (.A0(mult_29s_25s_0_pp_2_13), .A1(mult_29s_25s_0_pp_2_14), 
           .B0(mult_29s_25s_0_pp_3_13), .B1(mult_29s_25s_0_pp_3_14), .CI(co_mult_29s_25s_0_1_4), 
           .COUT(co_mult_29s_25s_0_1_5), .S0(s_mult_29s_25s_0_1_13), .S1(s_mult_29s_25s_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_6 (.A0(mult_29s_25s_0_pp_2_15), .A1(mult_29s_25s_0_pp_2_16), 
           .B0(mult_29s_25s_0_pp_3_15), .B1(mult_29s_25s_0_pp_3_16), .CI(co_mult_29s_25s_0_1_5), 
           .COUT(co_mult_29s_25s_0_1_6), .S0(s_mult_29s_25s_0_1_15), .S1(s_mult_29s_25s_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_7 (.A0(mult_29s_25s_0_pp_2_17), .A1(mult_29s_25s_0_pp_2_18), 
           .B0(mult_29s_25s_0_pp_3_17), .B1(mult_29s_25s_0_pp_3_18), .CI(co_mult_29s_25s_0_1_6), 
           .COUT(co_mult_29s_25s_0_1_7), .S0(s_mult_29s_25s_0_1_17), .S1(s_mult_29s_25s_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_8 (.A0(mult_29s_25s_0_pp_2_19), .A1(mult_29s_25s_0_pp_2_20), 
           .B0(mult_29s_25s_0_pp_3_19), .B1(mult_29s_25s_0_pp_3_20), .CI(co_mult_29s_25s_0_1_7), 
           .COUT(co_mult_29s_25s_0_1_8), .S0(s_mult_29s_25s_0_1_19), .S1(s_mult_29s_25s_0_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_9 (.A0(mult_29s_25s_0_pp_2_21), .A1(mult_29s_25s_0_pp_2_22), 
           .B0(mult_29s_25s_0_pp_3_21), .B1(mult_29s_25s_0_pp_3_22), .CI(co_mult_29s_25s_0_1_8), 
           .COUT(co_mult_29s_25s_0_1_9), .S0(s_mult_29s_25s_0_1_21), .S1(s_mult_29s_25s_0_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_10 (.A0(mult_29s_25s_0_pp_2_23), .A1(mult_29s_25s_0_pp_2_24), 
           .B0(mult_29s_25s_0_pp_3_23), .B1(mult_29s_25s_0_pp_3_24), .CI(co_mult_29s_25s_0_1_9), 
           .COUT(co_mult_29s_25s_0_1_10), .S0(s_mult_29s_25s_0_1_23), .S1(s_mult_29s_25s_0_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_11 (.A0(mult_29s_25s_0_pp_2_25), .A1(mult_29s_25s_0_pp_2_26), 
           .B0(mult_29s_25s_0_pp_3_25), .B1(mult_29s_25s_0_pp_3_26), .CI(co_mult_29s_25s_0_1_10), 
           .COUT(co_mult_29s_25s_0_1_11), .S0(s_mult_29s_25s_0_1_25), .S1(s_mult_29s_25s_0_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_1_12 (.A0(mult_29s_25s_0_pp_2_27), .A1(mult_29s_25s_0_pp_2_28), 
           .B0(mult_29s_25s_0_pp_3_27), .B1(mult_29s_25s_0_pp_3_28), .CI(co_mult_29s_25s_0_1_11), 
           .S0(s_mult_29s_25s_0_1_27), .S1(s_mult_29s_25s_0_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_2_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_4_10), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_5_10), .CI(GND_net), .COUT(co_mult_29s_25s_0_2_1), 
           .S1(s_mult_29s_25s_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_2 (.A0(mult_29s_25s_0_pp_4_11), .A1(mult_29s_25s_0_pp_4_12), 
           .B0(mult_29s_25s_0_pp_5_11), .B1(mult_29s_25s_0_pp_5_12), .CI(co_mult_29s_25s_0_2_1), 
           .COUT(co_mult_29s_25s_0_2_2), .S0(s_mult_29s_25s_0_2_11), .S1(s_mult_29s_25s_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_3 (.A0(mult_29s_25s_0_pp_4_13), .A1(mult_29s_25s_0_pp_4_14), 
           .B0(mult_29s_25s_0_pp_5_13), .B1(mult_29s_25s_0_pp_5_14), .CI(co_mult_29s_25s_0_2_2), 
           .COUT(co_mult_29s_25s_0_2_3), .S0(s_mult_29s_25s_0_2_13), .S1(s_mult_29s_25s_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_4 (.A0(mult_29s_25s_0_pp_4_15), .A1(mult_29s_25s_0_pp_4_16), 
           .B0(mult_29s_25s_0_pp_5_15), .B1(mult_29s_25s_0_pp_5_16), .CI(co_mult_29s_25s_0_2_3), 
           .COUT(co_mult_29s_25s_0_2_4), .S0(s_mult_29s_25s_0_2_15), .S1(s_mult_29s_25s_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_5 (.A0(mult_29s_25s_0_pp_4_17), .A1(mult_29s_25s_0_pp_4_18), 
           .B0(mult_29s_25s_0_pp_5_17), .B1(mult_29s_25s_0_pp_5_18), .CI(co_mult_29s_25s_0_2_4), 
           .COUT(co_mult_29s_25s_0_2_5), .S0(s_mult_29s_25s_0_2_17), .S1(s_mult_29s_25s_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_6 (.A0(mult_29s_25s_0_pp_4_19), .A1(mult_29s_25s_0_pp_4_20), 
           .B0(mult_29s_25s_0_pp_5_19), .B1(mult_29s_25s_0_pp_5_20), .CI(co_mult_29s_25s_0_2_5), 
           .COUT(co_mult_29s_25s_0_2_6), .S0(s_mult_29s_25s_0_2_19), .S1(s_mult_29s_25s_0_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_7 (.A0(mult_29s_25s_0_pp_4_21), .A1(mult_29s_25s_0_pp_4_22), 
           .B0(mult_29s_25s_0_pp_5_21), .B1(mult_29s_25s_0_pp_5_22), .CI(co_mult_29s_25s_0_2_6), 
           .COUT(co_mult_29s_25s_0_2_7), .S0(s_mult_29s_25s_0_2_21), .S1(s_mult_29s_25s_0_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_8 (.A0(mult_29s_25s_0_pp_4_23), .A1(mult_29s_25s_0_pp_4_24), 
           .B0(mult_29s_25s_0_pp_5_23), .B1(mult_29s_25s_0_pp_5_24), .CI(co_mult_29s_25s_0_2_7), 
           .COUT(co_mult_29s_25s_0_2_8), .S0(s_mult_29s_25s_0_2_23), .S1(s_mult_29s_25s_0_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_9 (.A0(mult_29s_25s_0_pp_4_25), .A1(mult_29s_25s_0_pp_4_26), 
           .B0(mult_29s_25s_0_pp_5_25), .B1(mult_29s_25s_0_pp_5_26), .CI(co_mult_29s_25s_0_2_8), 
           .COUT(co_mult_29s_25s_0_2_9), .S0(s_mult_29s_25s_0_2_25), .S1(s_mult_29s_25s_0_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_2_10 (.A0(mult_29s_25s_0_pp_4_27), .A1(mult_29s_25s_0_pp_4_28), 
           .B0(mult_29s_25s_0_pp_5_27), .B1(mult_29s_25s_0_pp_5_28), .CI(co_mult_29s_25s_0_2_9), 
           .S0(s_mult_29s_25s_0_2_27), .S1(s_mult_29s_25s_0_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_3_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_6_14), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_7_14), .CI(GND_net), .COUT(co_mult_29s_25s_0_3_1), 
           .S1(s_mult_29s_25s_0_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_2 (.A0(mult_29s_25s_0_pp_6_15), .A1(mult_29s_25s_0_pp_6_16), 
           .B0(mult_29s_25s_0_pp_7_15), .B1(mult_29s_25s_0_pp_7_16), .CI(co_mult_29s_25s_0_3_1), 
           .COUT(co_mult_29s_25s_0_3_2), .S0(s_mult_29s_25s_0_3_15), .S1(s_mult_29s_25s_0_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_3 (.A0(mult_29s_25s_0_pp_6_17), .A1(mult_29s_25s_0_pp_6_18), 
           .B0(mult_29s_25s_0_pp_7_17), .B1(mult_29s_25s_0_pp_7_18), .CI(co_mult_29s_25s_0_3_2), 
           .COUT(co_mult_29s_25s_0_3_3), .S0(s_mult_29s_25s_0_3_17), .S1(s_mult_29s_25s_0_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_4 (.A0(mult_29s_25s_0_pp_6_19), .A1(mult_29s_25s_0_pp_6_20), 
           .B0(mult_29s_25s_0_pp_7_19), .B1(mult_29s_25s_0_pp_7_20), .CI(co_mult_29s_25s_0_3_3), 
           .COUT(co_mult_29s_25s_0_3_4), .S0(s_mult_29s_25s_0_3_19), .S1(s_mult_29s_25s_0_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_5 (.A0(mult_29s_25s_0_pp_6_21), .A1(mult_29s_25s_0_pp_6_22), 
           .B0(mult_29s_25s_0_pp_7_21), .B1(mult_29s_25s_0_pp_7_22), .CI(co_mult_29s_25s_0_3_4), 
           .COUT(co_mult_29s_25s_0_3_5), .S0(s_mult_29s_25s_0_3_21), .S1(s_mult_29s_25s_0_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_6 (.A0(mult_29s_25s_0_pp_6_23), .A1(mult_29s_25s_0_pp_6_24), 
           .B0(mult_29s_25s_0_pp_7_23), .B1(mult_29s_25s_0_pp_7_24), .CI(co_mult_29s_25s_0_3_5), 
           .COUT(co_mult_29s_25s_0_3_6), .S0(s_mult_29s_25s_0_3_23), .S1(s_mult_29s_25s_0_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_7 (.A0(mult_29s_25s_0_pp_6_25), .A1(mult_29s_25s_0_pp_6_26), 
           .B0(mult_29s_25s_0_pp_7_25), .B1(mult_29s_25s_0_pp_7_26), .CI(co_mult_29s_25s_0_3_6), 
           .COUT(co_mult_29s_25s_0_3_7), .S0(s_mult_29s_25s_0_3_25), .S1(s_mult_29s_25s_0_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_3_8 (.A0(mult_29s_25s_0_pp_6_27), .A1(mult_29s_25s_0_pp_6_28), 
           .B0(mult_29s_25s_0_pp_7_27), .B1(mult_29s_25s_0_pp_7_28), .CI(co_mult_29s_25s_0_3_7), 
           .S0(s_mult_29s_25s_0_3_27), .S1(s_mult_29s_25s_0_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_4_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_8_18), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_9_18), .CI(GND_net), .COUT(co_mult_29s_25s_0_4_1), 
           .S1(s_mult_29s_25s_0_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_2 (.A0(mult_29s_25s_0_pp_8_19), .A1(mult_29s_25s_0_pp_8_20), 
           .B0(mult_29s_25s_0_pp_9_19), .B1(mult_29s_25s_0_pp_9_20), .CI(co_mult_29s_25s_0_4_1), 
           .COUT(co_mult_29s_25s_0_4_2), .S0(s_mult_29s_25s_0_4_19), .S1(s_mult_29s_25s_0_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_3 (.A0(mult_29s_25s_0_pp_8_21), .A1(mult_29s_25s_0_pp_8_22), 
           .B0(mult_29s_25s_0_pp_9_21), .B1(mult_29s_25s_0_pp_9_22), .CI(co_mult_29s_25s_0_4_2), 
           .COUT(co_mult_29s_25s_0_4_3), .S0(s_mult_29s_25s_0_4_21), .S1(s_mult_29s_25s_0_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_4 (.A0(mult_29s_25s_0_pp_8_23), .A1(mult_29s_25s_0_pp_8_24), 
           .B0(mult_29s_25s_0_pp_9_23), .B1(mult_29s_25s_0_pp_9_24), .CI(co_mult_29s_25s_0_4_3), 
           .COUT(co_mult_29s_25s_0_4_4), .S0(s_mult_29s_25s_0_4_23), .S1(s_mult_29s_25s_0_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_5 (.A0(mult_29s_25s_0_pp_8_25), .A1(mult_29s_25s_0_pp_8_26), 
           .B0(mult_29s_25s_0_pp_9_25), .B1(mult_29s_25s_0_pp_9_26), .CI(co_mult_29s_25s_0_4_4), 
           .COUT(co_mult_29s_25s_0_4_5), .S0(s_mult_29s_25s_0_4_25), .S1(s_mult_29s_25s_0_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_4_6 (.A0(mult_29s_25s_0_pp_8_27), .A1(mult_29s_25s_0_pp_8_28), 
           .B0(mult_29s_25s_0_pp_9_27), .B1(mult_29s_25s_0_pp_9_28), .CI(co_mult_29s_25s_0_4_5), 
           .S0(s_mult_29s_25s_0_4_27), .S1(s_mult_29s_25s_0_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_5_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_10_22), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_11_22), .CI(GND_net), .COUT(co_mult_29s_25s_0_5_1), 
           .S1(s_mult_29s_25s_0_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_2 (.A0(mult_29s_25s_0_pp_10_23), .A1(mult_29s_25s_0_pp_10_24), 
           .B0(mult_29s_25s_0_pp_11_23), .B1(mult_29s_25s_0_pp_11_24), .CI(co_mult_29s_25s_0_5_1), 
           .COUT(co_mult_29s_25s_0_5_2), .S0(s_mult_29s_25s_0_5_23), .S1(s_mult_29s_25s_0_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_3 (.A0(mult_29s_25s_0_pp_10_25), .A1(mult_29s_25s_0_pp_10_26), 
           .B0(mult_29s_25s_0_pp_11_25), .B1(mult_29s_25s_0_pp_11_26), .CI(co_mult_29s_25s_0_5_2), 
           .COUT(co_mult_29s_25s_0_5_3), .S0(s_mult_29s_25s_0_5_25), .S1(s_mult_29s_25s_0_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_5_4 (.A0(mult_29s_25s_0_pp_10_27), .A1(mult_29s_25s_0_pp_10_28), 
           .B0(mult_29s_25s_0_pp_11_27), .B1(mult_29s_25s_0_pp_11_28), .CI(co_mult_29s_25s_0_5_3), 
           .S0(s_mult_29s_25s_0_5_27), .S1(s_mult_29s_25s_0_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i13673_2_lut (.A(ss[3]), .B(ss[1]), .Z(n16258)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13673_2_lut.init = 16'heeee;
    FADD2B Cadd_mult_29s_25s_0_6_1 (.A0(GND_net), .A1(mult_29s_25s_0_pp_12_24), 
           .B0(GND_net), .B1(VCC_net), .CI(GND_net), .COUT(co_mult_29s_25s_0_6_1), 
           .S1(s_mult_29s_25s_0_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_2 (.A0(mult_29s_25s_0_pp_12_25), .A1(mult_29s_25s_0_pp_12_26), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_1), .COUT(co_mult_29s_25s_0_6_2), 
           .S0(s_mult_29s_25s_0_6_25), .S1(s_mult_29s_25s_0_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_6_3 (.A0(mult_29s_25s_0_pp_12_27), .A1(mult_29s_25s_0_pp_12_28), 
           .B0(GND_net), .B1(GND_net), .CI(co_mult_29s_25s_0_6_2), .S0(s_mult_29s_25s_0_6_27), 
           .S1(s_mult_29s_25s_0_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i3143_3_lut (.A(n3840), .B(n1068), .C(addOut[27]), .Z(intgOut0_28__N_1629[27])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3143_3_lut.init = 16'h3232;
    FADD2B Cadd_mult_29s_25s_0_7_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_0_4), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_2_4), .CI(GND_net), .COUT(co_mult_29s_25s_0_7_1), 
           .S1(multOut_28__N_1412[4])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_2 (.A0(s_mult_29s_25s_0_0_5), .A1(s_mult_29s_25s_0_0_6), 
           .B0(mult_29s_25s_0_pp_2_5), .B1(s_mult_29s_25s_0_1_6), .CI(co_mult_29s_25s_0_7_1), 
           .COUT(co_mult_29s_25s_0_7_2), .S0(multOut_28__N_1412[5]), .S1(multOut_28__N_1412[6])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_3 (.A0(s_mult_29s_25s_0_0_7), .A1(s_mult_29s_25s_0_0_8), 
           .B0(s_mult_29s_25s_0_1_7), .B1(s_mult_29s_25s_0_1_8), .CI(co_mult_29s_25s_0_7_2), 
           .COUT(co_mult_29s_25s_0_7_3), .S0(multOut_28__N_1412[7]), .S1(s_mult_29s_25s_0_7_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_4 (.A0(s_mult_29s_25s_0_0_9), .A1(s_mult_29s_25s_0_0_10), 
           .B0(s_mult_29s_25s_0_1_9), .B1(s_mult_29s_25s_0_1_10), .CI(co_mult_29s_25s_0_7_3), 
           .COUT(co_mult_29s_25s_0_7_4), .S0(s_mult_29s_25s_0_7_9), .S1(s_mult_29s_25s_0_7_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_5 (.A0(s_mult_29s_25s_0_0_11), .A1(s_mult_29s_25s_0_0_12), 
           .B0(s_mult_29s_25s_0_1_11), .B1(s_mult_29s_25s_0_1_12), .CI(co_mult_29s_25s_0_7_4), 
           .COUT(co_mult_29s_25s_0_7_5), .S0(s_mult_29s_25s_0_7_11), .S1(s_mult_29s_25s_0_7_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_6 (.A0(s_mult_29s_25s_0_0_13), .A1(s_mult_29s_25s_0_0_14), 
           .B0(s_mult_29s_25s_0_1_13), .B1(s_mult_29s_25s_0_1_14), .CI(co_mult_29s_25s_0_7_5), 
           .COUT(co_mult_29s_25s_0_7_6), .S0(s_mult_29s_25s_0_7_13), .S1(s_mult_29s_25s_0_7_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_7 (.A0(s_mult_29s_25s_0_0_15), .A1(s_mult_29s_25s_0_0_16), 
           .B0(s_mult_29s_25s_0_1_15), .B1(s_mult_29s_25s_0_1_16), .CI(co_mult_29s_25s_0_7_6), 
           .COUT(co_mult_29s_25s_0_7_7), .S0(s_mult_29s_25s_0_7_15), .S1(s_mult_29s_25s_0_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_8 (.A0(s_mult_29s_25s_0_0_17), .A1(s_mult_29s_25s_0_0_18), 
           .B0(s_mult_29s_25s_0_1_17), .B1(s_mult_29s_25s_0_1_18), .CI(co_mult_29s_25s_0_7_7), 
           .COUT(co_mult_29s_25s_0_7_8), .S0(s_mult_29s_25s_0_7_17), .S1(s_mult_29s_25s_0_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_9 (.A0(s_mult_29s_25s_0_0_19), .A1(s_mult_29s_25s_0_0_20), 
           .B0(s_mult_29s_25s_0_1_19), .B1(s_mult_29s_25s_0_1_20), .CI(co_mult_29s_25s_0_7_8), 
           .COUT(co_mult_29s_25s_0_7_9), .S0(s_mult_29s_25s_0_7_19), .S1(s_mult_29s_25s_0_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_10 (.A0(s_mult_29s_25s_0_0_21), .A1(s_mult_29s_25s_0_0_22), 
           .B0(s_mult_29s_25s_0_1_21), .B1(s_mult_29s_25s_0_1_22), .CI(co_mult_29s_25s_0_7_9), 
           .COUT(co_mult_29s_25s_0_7_10), .S0(s_mult_29s_25s_0_7_21), .S1(s_mult_29s_25s_0_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_11 (.A0(s_mult_29s_25s_0_0_23), .A1(s_mult_29s_25s_0_0_24), 
           .B0(s_mult_29s_25s_0_1_23), .B1(s_mult_29s_25s_0_1_24), .CI(co_mult_29s_25s_0_7_10), 
           .COUT(co_mult_29s_25s_0_7_11), .S0(s_mult_29s_25s_0_7_23), .S1(s_mult_29s_25s_0_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_12 (.A0(s_mult_29s_25s_0_0_25), .A1(s_mult_29s_25s_0_0_26), 
           .B0(s_mult_29s_25s_0_1_25), .B1(s_mult_29s_25s_0_1_26), .CI(co_mult_29s_25s_0_7_11), 
           .COUT(co_mult_29s_25s_0_7_12), .S0(s_mult_29s_25s_0_7_25), .S1(s_mult_29s_25s_0_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_7_13 (.A0(s_mult_29s_25s_0_0_27), .A1(s_mult_29s_25s_0_0_28), 
           .B0(s_mult_29s_25s_0_1_27), .B1(s_mult_29s_25s_0_1_28), .CI(co_mult_29s_25s_0_7_12), 
           .S0(s_mult_29s_25s_0_7_27), .S1(s_mult_29s_25s_0_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_8_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_2_12), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_6_12), .CI(GND_net), .COUT(co_mult_29s_25s_0_8_1), 
           .S1(s_mult_29s_25s_0_8_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_2 (.A0(s_mult_29s_25s_0_2_13), .A1(s_mult_29s_25s_0_2_14), 
           .B0(mult_29s_25s_0_pp_6_13), .B1(s_mult_29s_25s_0_3_14), .CI(co_mult_29s_25s_0_8_1), 
           .COUT(co_mult_29s_25s_0_8_2), .S0(s_mult_29s_25s_0_8_13), .S1(s_mult_29s_25s_0_8_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_3 (.A0(s_mult_29s_25s_0_2_15), .A1(s_mult_29s_25s_0_2_16), 
           .B0(s_mult_29s_25s_0_3_15), .B1(s_mult_29s_25s_0_3_16), .CI(co_mult_29s_25s_0_8_2), 
           .COUT(co_mult_29s_25s_0_8_3), .S0(s_mult_29s_25s_0_8_15), .S1(s_mult_29s_25s_0_8_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_4 (.A0(s_mult_29s_25s_0_2_17), .A1(s_mult_29s_25s_0_2_18), 
           .B0(s_mult_29s_25s_0_3_17), .B1(s_mult_29s_25s_0_3_18), .CI(co_mult_29s_25s_0_8_3), 
           .COUT(co_mult_29s_25s_0_8_4), .S0(s_mult_29s_25s_0_8_17), .S1(s_mult_29s_25s_0_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_5 (.A0(s_mult_29s_25s_0_2_19), .A1(s_mult_29s_25s_0_2_20), 
           .B0(s_mult_29s_25s_0_3_19), .B1(s_mult_29s_25s_0_3_20), .CI(co_mult_29s_25s_0_8_4), 
           .COUT(co_mult_29s_25s_0_8_5), .S0(s_mult_29s_25s_0_8_19), .S1(s_mult_29s_25s_0_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_6 (.A0(s_mult_29s_25s_0_2_21), .A1(s_mult_29s_25s_0_2_22), 
           .B0(s_mult_29s_25s_0_3_21), .B1(s_mult_29s_25s_0_3_22), .CI(co_mult_29s_25s_0_8_5), 
           .COUT(co_mult_29s_25s_0_8_6), .S0(s_mult_29s_25s_0_8_21), .S1(s_mult_29s_25s_0_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_7 (.A0(s_mult_29s_25s_0_2_23), .A1(s_mult_29s_25s_0_2_24), 
           .B0(s_mult_29s_25s_0_3_23), .B1(s_mult_29s_25s_0_3_24), .CI(co_mult_29s_25s_0_8_6), 
           .COUT(co_mult_29s_25s_0_8_7), .S0(s_mult_29s_25s_0_8_23), .S1(s_mult_29s_25s_0_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_8 (.A0(s_mult_29s_25s_0_2_25), .A1(s_mult_29s_25s_0_2_26), 
           .B0(s_mult_29s_25s_0_3_25), .B1(s_mult_29s_25s_0_3_26), .CI(co_mult_29s_25s_0_8_7), 
           .COUT(co_mult_29s_25s_0_8_8), .S0(s_mult_29s_25s_0_8_25), .S1(s_mult_29s_25s_0_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_8_9 (.A0(s_mult_29s_25s_0_2_27), .A1(s_mult_29s_25s_0_2_28), 
           .B0(s_mult_29s_25s_0_3_27), .B1(s_mult_29s_25s_0_3_28), .CI(co_mult_29s_25s_0_8_8), 
           .S0(s_mult_29s_25s_0_8_27), .S1(s_mult_29s_25s_0_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B Cadd_mult_29s_25s_0_9_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_4_20), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_10_20), .CI(GND_net), .COUT(co_mult_29s_25s_0_9_1), 
           .S1(s_mult_29s_25s_0_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_2 (.A0(s_mult_29s_25s_0_4_21), .A1(s_mult_29s_25s_0_4_22), 
           .B0(mult_29s_25s_0_pp_10_21), .B1(s_mult_29s_25s_0_5_22), .CI(co_mult_29s_25s_0_9_1), 
           .COUT(co_mult_29s_25s_0_9_2), .S0(s_mult_29s_25s_0_9_21), .S1(s_mult_29s_25s_0_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_3 (.A0(s_mult_29s_25s_0_4_23), .A1(s_mult_29s_25s_0_4_24), 
           .B0(s_mult_29s_25s_0_5_23), .B1(s_mult_29s_25s_0_5_24), .CI(co_mult_29s_25s_0_9_2), 
           .COUT(co_mult_29s_25s_0_9_3), .S0(s_mult_29s_25s_0_9_23), .S1(s_mult_29s_25s_0_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_4 (.A0(s_mult_29s_25s_0_4_25), .A1(s_mult_29s_25s_0_4_26), 
           .B0(s_mult_29s_25s_0_5_25), .B1(s_mult_29s_25s_0_5_26), .CI(co_mult_29s_25s_0_9_3), 
           .COUT(co_mult_29s_25s_0_9_4), .S0(s_mult_29s_25s_0_9_25), .S1(s_mult_29s_25s_0_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_9_5 (.A0(s_mult_29s_25s_0_4_27), .A1(s_mult_29s_25s_0_4_28), 
           .B0(s_mult_29s_25s_0_5_27), .B1(s_mult_29s_25s_0_5_28), .CI(co_mult_29s_25s_0_9_4), 
           .S0(s_mult_29s_25s_0_9_27), .S1(s_mult_29s_25s_0_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i19_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[18] ), 
         .D(\speed_avg_m2[18] ), .Z(subIn2_24__N_1348[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i18_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[17] ), 
         .D(\speed_avg_m2[17] ), .Z(subIn2_24__N_1348[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i18_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_mult_29s_25s_0_10_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_7_8), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_4_8), .CI(GND_net), .COUT(co_mult_29s_25s_0_10_1), 
           .S1(multOut_28__N_1412[8])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_2 (.A0(s_mult_29s_25s_0_7_9), .A1(s_mult_29s_25s_0_7_10), 
           .B0(mult_29s_25s_0_pp_4_9), .B1(s_mult_29s_25s_0_2_10), .CI(co_mult_29s_25s_0_10_1), 
           .COUT(co_mult_29s_25s_0_10_2), .S0(multOut_28__N_1412[9]), .S1(multOut_28__N_1412[10])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_3 (.A0(s_mult_29s_25s_0_7_11), .A1(s_mult_29s_25s_0_7_12), 
           .B0(s_mult_29s_25s_0_2_11), .B1(s_mult_29s_25s_0_8_12), .CI(co_mult_29s_25s_0_10_2), 
           .COUT(co_mult_29s_25s_0_10_3), .S0(multOut_28__N_1412[11]), .S1(multOut_28__N_1412[12])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_4 (.A0(s_mult_29s_25s_0_7_13), .A1(s_mult_29s_25s_0_7_14), 
           .B0(s_mult_29s_25s_0_8_13), .B1(s_mult_29s_25s_0_8_14), .CI(co_mult_29s_25s_0_10_3), 
           .COUT(co_mult_29s_25s_0_10_4), .S0(multOut_28__N_1412[13]), .S1(multOut_28__N_1412[14])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_5 (.A0(s_mult_29s_25s_0_7_15), .A1(s_mult_29s_25s_0_7_16), 
           .B0(s_mult_29s_25s_0_8_15), .B1(s_mult_29s_25s_0_8_16), .CI(co_mult_29s_25s_0_10_4), 
           .COUT(co_mult_29s_25s_0_10_5), .S0(multOut_28__N_1412[15]), .S1(s_mult_29s_25s_0_10_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_6 (.A0(s_mult_29s_25s_0_7_17), .A1(s_mult_29s_25s_0_7_18), 
           .B0(s_mult_29s_25s_0_8_17), .B1(s_mult_29s_25s_0_8_18), .CI(co_mult_29s_25s_0_10_5), 
           .COUT(co_mult_29s_25s_0_10_6), .S0(s_mult_29s_25s_0_10_17), .S1(s_mult_29s_25s_0_10_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_7 (.A0(s_mult_29s_25s_0_7_19), .A1(s_mult_29s_25s_0_7_20), 
           .B0(s_mult_29s_25s_0_8_19), .B1(s_mult_29s_25s_0_8_20), .CI(co_mult_29s_25s_0_10_6), 
           .COUT(co_mult_29s_25s_0_10_7), .S0(s_mult_29s_25s_0_10_19), .S1(s_mult_29s_25s_0_10_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_8 (.A0(s_mult_29s_25s_0_7_21), .A1(s_mult_29s_25s_0_7_22), 
           .B0(s_mult_29s_25s_0_8_21), .B1(s_mult_29s_25s_0_8_22), .CI(co_mult_29s_25s_0_10_7), 
           .COUT(co_mult_29s_25s_0_10_8), .S0(s_mult_29s_25s_0_10_21), .S1(s_mult_29s_25s_0_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_9 (.A0(s_mult_29s_25s_0_7_23), .A1(s_mult_29s_25s_0_7_24), 
           .B0(s_mult_29s_25s_0_8_23), .B1(s_mult_29s_25s_0_8_24), .CI(co_mult_29s_25s_0_10_8), 
           .COUT(co_mult_29s_25s_0_10_9), .S0(s_mult_29s_25s_0_10_23), .S1(s_mult_29s_25s_0_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_10 (.A0(s_mult_29s_25s_0_7_25), .A1(s_mult_29s_25s_0_7_26), 
           .B0(s_mult_29s_25s_0_8_25), .B1(s_mult_29s_25s_0_8_26), .CI(co_mult_29s_25s_0_10_9), 
           .COUT(co_mult_29s_25s_0_10_10), .S0(s_mult_29s_25s_0_10_25), 
           .S1(s_mult_29s_25s_0_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_10_11 (.A0(s_mult_29s_25s_0_7_27), .A1(s_mult_29s_25s_0_7_28), 
           .B0(s_mult_29s_25s_0_8_27), .B1(s_mult_29s_25s_0_8_28), .CI(co_mult_29s_25s_0_10_10), 
           .S0(s_mult_29s_25s_0_10_27), .S1(s_mult_29s_25s_0_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i17_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[16] ), 
         .D(\speed_avg_m2[16] ), .Z(subIn2_24__N_1348[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i17_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_223_15 (.A0(Out3[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18272), 
          .COUT(n18273), .S0(n1364[13]), .S1(n1364[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_15.INIT0 = 16'h5aaa;
    defparam add_223_15.INIT1 = 16'h5aaa;
    defparam add_223_15.INJECT1_0 = "NO";
    defparam add_223_15.INJECT1_1 = "NO";
    FADD2B Cadd_mult_29s_25s_0_11_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_9_24), 
           .B0(GND_net), .B1(s_mult_29s_25s_0_6_24), .CI(GND_net), .COUT(co_mult_29s_25s_0_11_1), 
           .S1(s_mult_29s_25s_0_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_2 (.A0(s_mult_29s_25s_0_9_25), .A1(s_mult_29s_25s_0_9_26), 
           .B0(s_mult_29s_25s_0_6_25), .B1(s_mult_29s_25s_0_6_26), .CI(co_mult_29s_25s_0_11_1), 
           .COUT(co_mult_29s_25s_0_11_2), .S0(s_mult_29s_25s_0_11_25), .S1(s_mult_29s_25s_0_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_add_11_3 (.A0(s_mult_29s_25s_0_9_27), .A1(s_mult_29s_25s_0_9_28), 
           .B0(s_mult_29s_25s_0_6_27), .B1(s_mult_29s_25s_0_6_28), .CI(co_mult_29s_25s_0_11_2), 
           .S0(s_mult_29s_25s_0_11_27), .S1(s_mult_29s_25s_0_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i16_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[15] ), 
         .D(\speed_avg_m2[15] ), .Z(subIn2_24__N_1348[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3368_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m2[2]), .Z(n5870)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3368_3_lut_4_lut.init = 16'hfd20;
    LUT4 subIn2_24__I_25_i15_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[14] ), 
         .D(\speed_avg_m2[14] ), .Z(subIn2_24__N_1348[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i15_3_lut_4_lut.init = 16'hfb40;
    FADD2B Cadd_t_mult_29s_25s_0_12_1 (.A0(GND_net), .A1(s_mult_29s_25s_0_10_16), 
           .B0(GND_net), .B1(mult_29s_25s_0_pp_8_16), .CI(GND_net), .COUT(co_t_mult_29s_25s_0_12_1), 
           .S1(multOut_28__N_1412[16])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_2 (.A0(s_mult_29s_25s_0_10_17), .A1(s_mult_29s_25s_0_10_18), 
           .B0(mult_29s_25s_0_pp_8_17), .B1(s_mult_29s_25s_0_4_18), .CI(co_t_mult_29s_25s_0_12_1), 
           .COUT(co_t_mult_29s_25s_0_12_2), .S0(multOut_28__N_1412[17]), 
           .S1(multOut_28__N_1412[18])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_3 (.A0(s_mult_29s_25s_0_10_19), .A1(s_mult_29s_25s_0_10_20), 
           .B0(s_mult_29s_25s_0_4_19), .B1(s_mult_29s_25s_0_9_20), .CI(co_t_mult_29s_25s_0_12_2), 
           .COUT(co_t_mult_29s_25s_0_12_3), .S0(multOut_28__N_1412[19]), 
           .S1(multOut_28__N_1412[20])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_4 (.A0(s_mult_29s_25s_0_10_21), .A1(s_mult_29s_25s_0_10_22), 
           .B0(s_mult_29s_25s_0_9_21), .B1(s_mult_29s_25s_0_9_22), .CI(co_t_mult_29s_25s_0_12_3), 
           .COUT(co_t_mult_29s_25s_0_12_4), .S0(multOut_28__N_1412[21]), 
           .S1(multOut_28__N_1412[22])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_5 (.A0(s_mult_29s_25s_0_10_23), .A1(s_mult_29s_25s_0_10_24), 
           .B0(s_mult_29s_25s_0_9_23), .B1(s_mult_29s_25s_0_11_24), .CI(co_t_mult_29s_25s_0_12_4), 
           .COUT(co_t_mult_29s_25s_0_12_5), .S0(multOut_28__N_1412[23]), 
           .S1(multOut_28__N_1412[24])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_6 (.A0(s_mult_29s_25s_0_10_25), .A1(s_mult_29s_25s_0_10_26), 
           .B0(s_mult_29s_25s_0_11_25), .B1(s_mult_29s_25s_0_11_26), .CI(co_t_mult_29s_25s_0_12_5), 
           .COUT(co_t_mult_29s_25s_0_12_6), .S0(multOut_28__N_1412[25]), 
           .S1(multOut_28__N_1412[26])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B t_mult_29s_25s_0_add_12_7 (.A0(s_mult_29s_25s_0_10_27), .A1(s_mult_29s_25s_0_10_28), 
           .B0(s_mult_29s_25s_0_11_27), .B1(s_mult_29s_25s_0_11_28), .CI(co_t_mult_29s_25s_0_12_6), 
           .S0(multOut_28__N_1412[27]), .S1(multOut_28__N_1412[28])) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i3141_3_lut (.A(n3840), .B(n1068), .C(addOut[26]), .Z(intgOut0_28__N_1629[26])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3141_3_lut.init = 16'h3232;
    MULT2 mult_29s_25s_0_mult_0_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mult_29s_25s_0_cin_lr_0), .CO(mco), .P0(multOut_28__N_1412[1]), 
          .P1(mult_29s_25s_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco), .CO(mco_1), .P0(mult_29s_25s_0_pp_0_3), 
          .P1(mult_29s_25s_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_1), .CO(mco_2), .P0(mult_29s_25s_0_pp_0_5), 
          .P1(mult_29s_25s_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_2), .CO(mco_3), .P0(mult_29s_25s_0_pp_0_7), 
          .P1(mult_29s_25s_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_3), .CO(mco_4), .P0(mult_29s_25s_0_pp_0_9), 
          .P1(mult_29s_25s_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_4), .CO(mco_5), .P0(mult_29s_25s_0_pp_0_11), 
          .P1(mult_29s_25s_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_5), .CO(mco_6), .P0(mult_29s_25s_0_pp_0_13), 
          .P1(mult_29s_25s_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_6), .CO(mco_7), .P0(mult_29s_25s_0_pp_0_15), 
          .P1(mult_29s_25s_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_7), .CO(mco_8), .P0(mult_29s_25s_0_pp_0_17), 
          .P1(mult_29s_25s_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_8), .CO(mco_9), .P0(mult_29s_25s_0_pp_0_19), 
          .P1(mult_29s_25s_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_9), .CO(mco_10), .P0(mult_29s_25s_0_pp_0_21), 
          .P1(mult_29s_25s_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_10), .CO(mco_11), .P0(mult_29s_25s_0_pp_0_23), 
          .P1(mult_29s_25s_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_11), .CO(mco_12), .P0(mult_29s_25s_0_pp_0_25), 
          .P1(mult_29s_25s_0_pp_0_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_0_13 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(GND_net), .B1(multIn2[0]), .B2(GND_net), 
          .B3(multIn2[0]), .CI(mco_12), .P0(mult_29s_25s_0_pp_0_27), .P1(mult_29s_25s_0_pp_0_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_2), .CO(mco_14), .P0(mult_29s_25s_0_pp_1_3), 
          .P1(mult_29s_25s_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_14), .CO(mco_15), .P0(mult_29s_25s_0_pp_1_5), 
          .P1(mult_29s_25s_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_15), .CO(mco_16), .P0(mult_29s_25s_0_pp_1_7), 
          .P1(mult_29s_25s_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_16), .CO(mco_17), .P0(mult_29s_25s_0_pp_1_9), 
          .P1(mult_29s_25s_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_17), .CO(mco_18), .P0(mult_29s_25s_0_pp_1_11), 
          .P1(mult_29s_25s_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_18), .CO(mco_19), .P0(mult_29s_25s_0_pp_1_13), 
          .P1(mult_29s_25s_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_19), .CO(mco_20), .P0(mult_29s_25s_0_pp_1_15), 
          .P1(mult_29s_25s_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_20), .CO(mco_21), .P0(mult_29s_25s_0_pp_1_17), 
          .P1(mult_29s_25s_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_21), .CO(mco_22), .P0(mult_29s_25s_0_pp_1_19), 
          .P1(mult_29s_25s_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_22), .CO(mco_23), .P0(mult_29s_25s_0_pp_1_21), 
          .P1(mult_29s_25s_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_23), .CO(mco_24), .P0(mult_29s_25s_0_pp_1_23), 
          .P1(mult_29s_25s_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_24), .CO(mco_25), .P0(mult_29s_25s_0_pp_1_25), 
          .P1(mult_29s_25s_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_2_12 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[3]), .B1(GND_net), .B2(multIn2[3]), 
          .B3(GND_net), .CI(mco_25), .P0(mult_29s_25s_0_pp_1_27), .P1(mult_29s_25s_0_pp_1_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_4), .CO(mco_28), .P0(mult_29s_25s_0_pp_2_5), 
          .P1(mult_29s_25s_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_28), .CO(mco_29), .P0(mult_29s_25s_0_pp_2_7), 
          .P1(mult_29s_25s_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_29), .CO(mco_30), .P0(mult_29s_25s_0_pp_2_9), 
          .P1(mult_29s_25s_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_30), .CO(mco_31), .P0(mult_29s_25s_0_pp_2_11), 
          .P1(mult_29s_25s_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_31), .CO(mco_32), .P0(mult_29s_25s_0_pp_2_13), 
          .P1(mult_29s_25s_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_32), .CO(mco_33), .P0(mult_29s_25s_0_pp_2_15), 
          .P1(mult_29s_25s_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_33), .CO(mco_34), .P0(mult_29s_25s_0_pp_2_17), 
          .P1(mult_29s_25s_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_34), .CO(mco_35), .P0(mult_29s_25s_0_pp_2_19), 
          .P1(mult_29s_25s_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_35), .CO(mco_36), .P0(mult_29s_25s_0_pp_2_21), 
          .P1(mult_29s_25s_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_36), .CO(mco_37), .P0(mult_29s_25s_0_pp_2_23), 
          .P1(mult_29s_25s_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_37), .CO(mco_38), .P0(mult_29s_25s_0_pp_2_25), 
          .P1(mult_29s_25s_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_4_11 (.A0(subOut[23]), .A1(subOut[23]), .A2(subOut[23]), 
          .A3(subOut[23]), .B0(multIn2[9]), .B1(GND_net), .B2(multIn2[9]), 
          .B3(GND_net), .CI(mco_38), .P0(mult_29s_25s_0_pp_2_27), .P1(mult_29s_25s_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i14_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[13] ), 
         .D(\speed_avg_m2[13] ), .Z(subIn2_24__N_1348[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i14_3_lut_4_lut.init = 16'hfb40;
    MULT2 mult_29s_25s_0_mult_6_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mult_29s_25s_0_cin_lr_6), .CO(mco_42), 
          .P0(mult_29s_25s_0_pp_3_7), .P1(mult_29s_25s_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_42), .CO(mco_43), .P0(mult_29s_25s_0_pp_3_9), 
          .P1(mult_29s_25s_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_43), .CO(mco_44), .P0(mult_29s_25s_0_pp_3_11), 
          .P1(mult_29s_25s_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_44), .CO(mco_45), .P0(mult_29s_25s_0_pp_3_13), 
          .P1(mult_29s_25s_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_45), .CO(mco_46), .P0(mult_29s_25s_0_pp_3_15), 
          .P1(mult_29s_25s_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_46), .CO(mco_47), .P0(mult_29s_25s_0_pp_3_17), 
          .P1(mult_29s_25s_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_47), .CO(mco_48), .P0(mult_29s_25s_0_pp_3_19), 
          .P1(mult_29s_25s_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_48), .CO(mco_49), .P0(mult_29s_25s_0_pp_3_21), 
          .P1(mult_29s_25s_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_49), .CO(mco_50), .P0(mult_29s_25s_0_pp_3_23), 
          .P1(mult_29s_25s_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_50), .CO(mco_51), .P0(mult_29s_25s_0_pp_3_25), 
          .P1(mult_29s_25s_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_6_10 (.A0(subOut[20]), .A1(subOut[21]), .A2(subOut[21]), 
          .A3(subOut[23]), .B0(multIn2[9]), .B1(multIn2[3]), .B2(multIn2[9]), 
          .B3(multIn2[3]), .CI(mco_51), .P0(mult_29s_25s_0_pp_3_27), .P1(mult_29s_25s_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mult_29s_25s_0_cin_lr_8), .CO(mco_56), 
          .P0(mult_29s_25s_0_pp_4_9), .P1(mult_29s_25s_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_56), .CO(mco_57), .P0(mult_29s_25s_0_pp_4_11), 
          .P1(mult_29s_25s_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_57), .CO(mco_58), .P0(mult_29s_25s_0_pp_4_13), 
          .P1(mult_29s_25s_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_58), .CO(mco_59), .P0(mult_29s_25s_0_pp_4_15), 
          .P1(mult_29s_25s_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_59), .CO(mco_60), .P0(mult_29s_25s_0_pp_4_17), 
          .P1(mult_29s_25s_0_pp_4_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_60), .CO(mco_61), .P0(mult_29s_25s_0_pp_4_19), 
          .P1(mult_29s_25s_0_pp_4_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_61), .CO(mco_62), .P0(mult_29s_25s_0_pp_4_21), 
          .P1(mult_29s_25s_0_pp_4_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_62), .CO(mco_63), .P0(mult_29s_25s_0_pp_4_23), 
          .P1(mult_29s_25s_0_pp_4_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_63), .CO(mco_64), .P0(mult_29s_25s_0_pp_4_25), 
          .P1(mult_29s_25s_0_pp_4_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_8_9 (.A0(subOut[18]), .A1(subOut[19]), .A2(subOut[19]), 
          .A3(subOut[20]), .B0(multIn2[9]), .B1(multIn2[9]), .B2(multIn2[9]), 
          .B3(multIn2[9]), .CI(mco_64), .P0(mult_29s_25s_0_pp_4_27), .P1(mult_29s_25s_0_pp_4_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mult_29s_25s_0_cin_lr_10), .CO(mco_70), 
          .P0(mult_29s_25s_0_pp_5_11), .P1(mult_29s_25s_0_pp_5_12)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_70), .CO(mco_71), .P0(mult_29s_25s_0_pp_5_13), 
          .P1(mult_29s_25s_0_pp_5_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_71), .CO(mco_72), .P0(mult_29s_25s_0_pp_5_15), 
          .P1(mult_29s_25s_0_pp_5_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_72), .CO(mco_73), .P0(mult_29s_25s_0_pp_5_17), 
          .P1(mult_29s_25s_0_pp_5_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_73), .CO(mco_74), .P0(mult_29s_25s_0_pp_5_19), 
          .P1(mult_29s_25s_0_pp_5_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_74), .CO(mco_75), .P0(mult_29s_25s_0_pp_5_21), 
          .P1(mult_29s_25s_0_pp_5_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_75), .CO(mco_76), .P0(mult_29s_25s_0_pp_5_23), 
          .P1(mult_29s_25s_0_pp_5_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_76), .CO(mco_77), .P0(mult_29s_25s_0_pp_5_25), 
          .P1(mult_29s_25s_0_pp_5_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_10_8 (.A0(subOut[16]), .A1(subOut[17]), .A2(subOut[17]), 
          .A3(subOut[18]), .B0(multIn2[11]), .B1(multIn2[11]), .B2(multIn2[11]), 
          .B3(multIn2[11]), .CI(mco_77), .P0(mult_29s_25s_0_pp_5_27), 
          .P1(mult_29s_25s_0_pp_5_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i12_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[11] ), 
         .D(\speed_avg_m2[11] ), .Z(subIn2_24__N_1348[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i12_3_lut_4_lut.init = 16'hfb40;
    MULT2 mult_29s_25s_0_mult_12_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_12), .CO(mco_84), .P0(mult_29s_25s_0_pp_6_13), 
          .P1(mult_29s_25s_0_pp_6_14)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_84), .CO(mco_85), .P0(mult_29s_25s_0_pp_6_15), 
          .P1(mult_29s_25s_0_pp_6_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_85), .CO(mco_86), .P0(mult_29s_25s_0_pp_6_17), 
          .P1(mult_29s_25s_0_pp_6_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_86), .CO(mco_87), .P0(mult_29s_25s_0_pp_6_19), 
          .P1(mult_29s_25s_0_pp_6_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_87), .CO(mco_88), .P0(mult_29s_25s_0_pp_6_21), 
          .P1(mult_29s_25s_0_pp_6_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_88), .CO(mco_89), .P0(mult_29s_25s_0_pp_6_23), 
          .P1(mult_29s_25s_0_pp_6_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_89), .CO(mco_90), .P0(mult_29s_25s_0_pp_6_25), 
          .P1(mult_29s_25s_0_pp_6_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_12_7 (.A0(subOut[14]), .A1(subOut[15]), .A2(subOut[15]), 
          .A3(subOut[16]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_90), .P0(mult_29s_25s_0_pp_6_27), .P1(mult_29s_25s_0_pp_6_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_14), .CO(mco_98), .P0(mult_29s_25s_0_pp_7_15), 
          .P1(mult_29s_25s_0_pp_7_16)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_98), .CO(mco_99), .P0(mult_29s_25s_0_pp_7_17), 
          .P1(mult_29s_25s_0_pp_7_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_99), .CO(mco_100), .P0(mult_29s_25s_0_pp_7_19), 
          .P1(mult_29s_25s_0_pp_7_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_100), .CO(mco_101), .P0(mult_29s_25s_0_pp_7_21), 
          .P1(mult_29s_25s_0_pp_7_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_101), .CO(mco_102), .P0(mult_29s_25s_0_pp_7_23), 
          .P1(mult_29s_25s_0_pp_7_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_102), .CO(mco_103), .P0(mult_29s_25s_0_pp_7_25), 
          .P1(mult_29s_25s_0_pp_7_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_14_6 (.A0(subOut[12]), .A1(subOut[13]), .A2(subOut[13]), 
          .A3(subOut[14]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_103), .P0(mult_29s_25s_0_pp_7_27), .P1(mult_29s_25s_0_pp_7_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_16), .CO(mco_112), .P0(mult_29s_25s_0_pp_8_17), 
          .P1(mult_29s_25s_0_pp_8_18)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_112), .CO(mco_113), .P0(mult_29s_25s_0_pp_8_19), 
          .P1(mult_29s_25s_0_pp_8_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_113), .CO(mco_114), .P0(mult_29s_25s_0_pp_8_21), 
          .P1(mult_29s_25s_0_pp_8_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_114), .CO(mco_115), .P0(mult_29s_25s_0_pp_8_23), 
          .P1(mult_29s_25s_0_pp_8_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_115), .CO(mco_116), .P0(mult_29s_25s_0_pp_8_25), 
          .P1(mult_29s_25s_0_pp_8_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_16_5 (.A0(subOut[10]), .A1(subOut[11]), .A2(subOut[11]), 
          .A3(subOut[12]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_116), .P0(mult_29s_25s_0_pp_8_27), .P1(mult_29s_25s_0_pp_8_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_18), .CO(mco_126), .P0(mult_29s_25s_0_pp_9_19), 
          .P1(mult_29s_25s_0_pp_9_20)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_126), .CO(mco_127), .P0(mult_29s_25s_0_pp_9_21), 
          .P1(mult_29s_25s_0_pp_9_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_127), .CO(mco_128), .P0(mult_29s_25s_0_pp_9_23), 
          .P1(mult_29s_25s_0_pp_9_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_128), .CO(mco_129), .P0(mult_29s_25s_0_pp_9_25), 
          .P1(mult_29s_25s_0_pp_9_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_18_4 (.A0(subOut[8]), .A1(subOut[9]), .A2(subOut[9]), 
          .A3(subOut[10]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_129), .P0(mult_29s_25s_0_pp_9_27), .P1(mult_29s_25s_0_pp_9_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 i3139_3_lut (.A(n3840), .B(n1068), .C(addOut[25]), .Z(intgOut0_28__N_1629[25])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3139_3_lut.init = 16'h3232;
    MULT2 mult_29s_25s_0_mult_20_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_20), .CO(mco_140), .P0(mult_29s_25s_0_pp_10_21), 
          .P1(mult_29s_25s_0_pp_10_22)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_140), .CO(mco_141), .P0(mult_29s_25s_0_pp_10_23), 
          .P1(mult_29s_25s_0_pp_10_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_141), .CO(mco_142), .P0(mult_29s_25s_0_pp_10_25), 
          .P1(mult_29s_25s_0_pp_10_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_20_3 (.A0(subOut[6]), .A1(subOut[7]), .A2(subOut[7]), 
          .A3(subOut[8]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_142), .P0(mult_29s_25s_0_pp_10_27), .P1(mult_29s_25s_0_pp_10_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_0 (.A0(subOut[0]), .A1(subOut[1]), .A2(subOut[1]), 
          .A3(subOut[2]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mult_29s_25s_0_cin_lr_22), .CO(mco_154), .P0(mult_29s_25s_0_pp_11_23), 
          .P1(mult_29s_25s_0_pp_11_24)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_1 (.A0(subOut[2]), .A1(subOut[3]), .A2(subOut[3]), 
          .A3(subOut[4]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_154), .CO(mco_155), .P0(mult_29s_25s_0_pp_11_25), 
          .P1(mult_29s_25s_0_pp_11_26)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    MULT2 mult_29s_25s_0_mult_22_2 (.A0(subOut[4]), .A1(subOut[5]), .A2(subOut[5]), 
          .A3(subOut[6]), .B0(GND_net), .B1(GND_net), .B2(GND_net), 
          .B3(GND_net), .CI(mco_155), .P0(mult_29s_25s_0_pp_11_27), .P1(mult_29s_25s_0_pp_11_28)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    FADD2B mult_29s_25s_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_29s_25s_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(229[14:21])
    LUT4 subIn2_24__I_25_i11_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[10] ), 
         .D(\speed_avg_m2[10] ), .Z(subIn2_24__N_1348[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i7_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[6] ), 
         .D(\speed_avg_m2[6] ), .Z(subIn2_24__N_1348[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i6_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[5] ), 
         .D(\speed_avg_m2[5] ), .Z(subIn2_24__N_1348[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i5_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[4] ), 
         .D(\speed_avg_m2[4] ), .Z(subIn2_24__N_1348[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 ss_4__I_0_353_i6_2_lut (.A(ss[0]), .B(ss[1]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(165[9:16])
    defparam ss_4__I_0_353_i6_2_lut.init = 16'heeee;
    LUT4 subIn2_24__I_25_i3_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[2] ), 
         .D(\speed_avg_m2[2] ), .Z(subIn2_24__N_1348[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13250_2_lut (.A(addOut[0]), .B(n22216), .Z(Out3_28__N_1174[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13250_2_lut.init = 16'h2222;
    LUT4 mux_92_i10_3_lut (.A(\speed_avg_m3[9] ), .B(\speed_avg_m2[9] ), 
         .C(n22204), .Z(subIn2_24__N_1535[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i10_3_lut.init = 16'hcaca;
    LUT4 subIn2_24__I_25_i2_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[1] ), 
         .D(\speed_avg_m2[1] ), .Z(subIn2_24__N_1348[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 subIn2_24__I_25_i1_3_lut_4_lut (.A(ss[2]), .B(n21470), .C(\speed_avg_m1[0] ), 
         .D(\speed_avg_m2[0] ), .Z(subIn2_24__N_1348[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam subIn2_24__I_25_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_3_lut_4_lut (.A(ss[3]), .B(n21492), .C(ss[0]), .D(n22216), 
         .Z(multIn2[11])) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(96[9:11])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0060;
    LUT4 i3370_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m2[3]), .Z(n5872)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3370_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3137_3_lut (.A(n3840), .B(n1068), .C(addOut[24]), .Z(intgOut0_28__N_1629[24])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3137_3_lut.init = 16'h3232;
    LUT4 i1_4_lut_adj_59 (.A(n21498), .B(ss[3]), .C(ss[0]), .D(ss[1]), 
         .Z(subIn1_24__N_1342)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_adj_59.init = 16'h0150;
    LUT4 i2_4_lut_adj_60 (.A(n21409), .B(n15757), .C(n21408), .D(n56), 
         .Z(n16223)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i2_4_lut_adj_60.init = 16'hfbfa;
    LUT4 i3135_3_lut (.A(n3840), .B(n1068), .C(addOut[23]), .Z(intgOut0_28__N_1629[23])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3135_3_lut.init = 16'h3232;
    LUT4 i1_3_lut_4_lut (.A(n1068), .B(n3840), .C(n21427), .D(clk_N_875_enable_392), 
         .Z(n15143)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfe00;
    LUT4 i1_4_lut_4_lut_adj_61 (.A(n21403), .B(n16223), .C(n21404), .D(n21405), 
         .Z(n19649)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam i1_4_lut_4_lut_adj_61.init = 16'h5400;
    LUT4 i3133_3_lut (.A(n3840), .B(n1068), .C(addOut[22]), .Z(intgOut0_28__N_1629[22])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3133_3_lut.init = 16'h3232;
    LUT4 i3372_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m2[4]), .Z(n5874)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3372_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX backOut0_i0_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut0_i0_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_69), 
            .CK(clk_N_875), .Q(backOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut0_i0_i1.GSR = "DISABLED";
    FD1S3AX multOut_i1 (.D(multOut_28__N_1412[1]), .CK(clk_N_875), .Q(multOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i1.GSR = "ENABLED";
    LUT4 mux_92_i9_3_lut (.A(\speed_avg_m3[8] ), .B(\speed_avg_m2[8] ), 
         .C(n22204), .Z(subIn2_24__N_1535[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i9_3_lut.init = 16'hcaca;
    LUT4 i11570_3_lut_4_lut (.A(n1068), .B(n3840), .C(n21438), .D(clk_N_875_enable_387), 
         .Z(n14299)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i11570_3_lut_4_lut.init = 16'hfe00;
    LUT4 i3374_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m2[5]), .Z(n5876)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3374_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i8_3_lut (.A(\speed_avg_m3[7] ), .B(\speed_avg_m2[7] ), 
         .C(n22204), .Z(subIn2_24__N_1535[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i8_3_lut.init = 16'hcaca;
    LUT4 i3131_3_lut (.A(n3840), .B(n1068), .C(addOut[20]), .Z(intgOut0_28__N_1629[20])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3131_3_lut.init = 16'h3232;
    LUT4 i3129_3_lut (.A(n3840), .B(n1068), .C(addOut[17]), .Z(intgOut0_28__N_1629[17])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3129_3_lut.init = 16'h3232;
    LUT4 mux_92_i4_3_lut (.A(\speed_avg_m3[3] ), .B(\speed_avg_m2[3] ), 
         .C(n22204), .Z(subIn2_24__N_1535[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i4_3_lut.init = 16'hcaca;
    LUT4 mux_92_i20_4_lut (.A(\speed_avg_m4[19] ), .B(\speed_avg_m3[19] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i20_4_lut.init = 16'hcac0;
    LUT4 i7_4_lut (.A(Out3[3]), .B(n14_adj_2334), .C(n10_adj_2335), .D(Out3[4]), 
         .Z(n18754)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut (.A(Out3[11]), .B(Out3[7]), .C(Out3[2]), .D(Out3[10]), 
         .Z(n14_adj_2334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_adj_62 (.A(Out3[9]), .B(Out3[1]), .Z(n10_adj_2335)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i2_2_lut_adj_62.init = 16'heeee;
    LUT4 i4_4_lut_adj_63 (.A(Out3[5]), .B(Out3[6]), .C(Out3[0]), .D(n6_adj_2336), 
         .Z(n18755)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i4_4_lut_adj_63.init = 16'hfffe;
    LUT4 i3127_3_lut (.A(n3840), .B(n1068), .C(addOut[13]), .Z(intgOut0_28__N_1629[13])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3127_3_lut.init = 16'h3232;
    LUT4 mux_92_i19_4_lut (.A(\speed_avg_m4[18] ), .B(\speed_avg_m3[18] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i19_4_lut.init = 16'hcac0;
    LUT4 i3376_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m2[6]), .Z(n5878)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3376_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3378_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[7]), 
         .D(speed_set_m2[7]), .Z(n5880)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3378_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_64 (.A(ss[3]), .B(n19662), .C(n22216), .D(n21462), 
         .Z(clk_N_875_enable_41)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_64.init = 16'hc4c0;
    LUT4 i3125_3_lut (.A(n3840), .B(n1068), .C(addOut[12]), .Z(intgOut0_28__N_1629[12])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3125_3_lut.init = 16'h3232;
    LUT4 i1_2_lut (.A(Out3[8]), .B(Out3[12]), .Z(n6_adj_2336)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i3123_3_lut (.A(n3840), .B(n1068), .C(addOut[11]), .Z(intgOut0_28__N_1629[11])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3123_3_lut.init = 16'h3232;
    LUT4 i7_4_lut_adj_65 (.A(Out2[3]), .B(n14_adj_2337), .C(n10_adj_2338), 
         .D(Out2[4]), .Z(n18757)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i7_4_lut_adj_65.init = 16'hfffe;
    LUT4 mux_92_i18_4_lut (.A(\speed_avg_m4[17] ), .B(\speed_avg_m3[17] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i18_4_lut.init = 16'hcac0;
    LUT4 i3121_3_lut (.A(n3840), .B(n1068), .C(addOut[8]), .Z(intgOut0_28__N_1629[8])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(267[4] 273[11])
    defparam i3121_3_lut.init = 16'h3232;
    LUT4 i6_4_lut_adj_66 (.A(Out2[11]), .B(Out2[7]), .C(Out2[2]), .D(Out2[10]), 
         .Z(n14_adj_2337)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i6_4_lut_adj_66.init = 16'hfffe;
    LUT4 mux_92_i17_4_lut (.A(\speed_avg_m4[16] ), .B(\speed_avg_m3[16] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i17_4_lut.init = 16'hcac0;
    LUT4 mux_92_i16_4_lut (.A(\speed_avg_m4[15] ), .B(\speed_avg_m3[15] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i16_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_rep_303 (.A(subIn1_24__N_1342), .B(n35), .Z(n21404)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam i1_2_lut_rep_303.init = 16'h8888;
    LUT4 i2_2_lut_adj_67 (.A(Out2[9]), .B(Out2[1]), .Z(n10_adj_2338)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i2_2_lut_adj_67.init = 16'heeee;
    LUT4 i1_4_lut_adj_68 (.A(n21492), .B(n19662), .C(n22216), .D(n11644), 
         .Z(clk_N_875_enable_209)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_68.init = 16'hc4c0;
    LUT4 i4_4_lut_adj_69 (.A(Out2[5]), .B(Out2[6]), .C(Out2[0]), .D(n6_adj_2339), 
         .Z(n18758)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i4_4_lut_adj_69.init = 16'hfffe;
    FD1S3AX multOut_i2 (.D(multOut_28__N_1412[2]), .CK(clk_N_875), .Q(multOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i2.GSR = "ENABLED";
    FD1S3AX multOut_i3 (.D(multOut_28__N_1412[3]), .CK(clk_N_875), .Q(multOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i3.GSR = "ENABLED";
    FD1S3AX multOut_i4 (.D(multOut_28__N_1412[4]), .CK(clk_N_875), .Q(multOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i4.GSR = "ENABLED";
    FD1S3AX multOut_i5 (.D(multOut_28__N_1412[5]), .CK(clk_N_875), .Q(multOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i5.GSR = "ENABLED";
    FD1S3AX multOut_i6 (.D(multOut_28__N_1412[6]), .CK(clk_N_875), .Q(multOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i6.GSR = "ENABLED";
    FD1S3AX multOut_i7 (.D(multOut_28__N_1412[7]), .CK(clk_N_875), .Q(multOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i7.GSR = "ENABLED";
    FD1S3AX multOut_i8 (.D(multOut_28__N_1412[8]), .CK(clk_N_875), .Q(multOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i8.GSR = "ENABLED";
    FD1S3AX multOut_i9 (.D(multOut_28__N_1412[9]), .CK(clk_N_875), .Q(multOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i9.GSR = "ENABLED";
    FD1S3AX multOut_i10 (.D(multOut_28__N_1412[10]), .CK(clk_N_875), .Q(multOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i10.GSR = "ENABLED";
    FD1S3AX multOut_i11 (.D(multOut_28__N_1412[11]), .CK(clk_N_875), .Q(multOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i11.GSR = "ENABLED";
    FD1S3AX multOut_i12 (.D(multOut_28__N_1412[12]), .CK(clk_N_875), .Q(multOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i12.GSR = "ENABLED";
    FD1S3AX multOut_i13 (.D(multOut_28__N_1412[13]), .CK(clk_N_875), .Q(multOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i13.GSR = "ENABLED";
    FD1S3AX multOut_i14 (.D(multOut_28__N_1412[14]), .CK(clk_N_875), .Q(multOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i14.GSR = "ENABLED";
    FD1S3AX multOut_i15 (.D(multOut_28__N_1412[15]), .CK(clk_N_875), .Q(multOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i15.GSR = "ENABLED";
    FD1S3AX multOut_i16 (.D(multOut_28__N_1412[16]), .CK(clk_N_875), .Q(multOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i16.GSR = "ENABLED";
    FD1S3AX multOut_i17 (.D(multOut_28__N_1412[17]), .CK(clk_N_875), .Q(multOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i17.GSR = "ENABLED";
    FD1S3AX multOut_i18 (.D(multOut_28__N_1412[18]), .CK(clk_N_875), .Q(multOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i18.GSR = "ENABLED";
    FD1S3AX multOut_i19 (.D(multOut_28__N_1412[19]), .CK(clk_N_875), .Q(multOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i19.GSR = "ENABLED";
    FD1S3AX multOut_i20 (.D(multOut_28__N_1412[20]), .CK(clk_N_875), .Q(multOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i20.GSR = "ENABLED";
    FD1S3AX multOut_i21 (.D(multOut_28__N_1412[21]), .CK(clk_N_875), .Q(multOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i21.GSR = "ENABLED";
    FD1S3AX multOut_i22 (.D(multOut_28__N_1412[22]), .CK(clk_N_875), .Q(multOut[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i22.GSR = "ENABLED";
    FD1S3AX multOut_i23 (.D(multOut_28__N_1412[23]), .CK(clk_N_875), .Q(multOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i23.GSR = "ENABLED";
    FD1S3AX multOut_i24 (.D(multOut_28__N_1412[24]), .CK(clk_N_875), .Q(multOut[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i24.GSR = "ENABLED";
    FD1S3AX multOut_i25 (.D(multOut_28__N_1412[25]), .CK(clk_N_875), .Q(multOut[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i25.GSR = "ENABLED";
    FD1S3AX multOut_i26 (.D(multOut_28__N_1412[26]), .CK(clk_N_875), .Q(multOut[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i26.GSR = "ENABLED";
    FD1S3AX multOut_i27 (.D(multOut_28__N_1412[27]), .CK(clk_N_875), .Q(multOut[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i27.GSR = "ENABLED";
    FD1S3AX multOut_i28 (.D(multOut_28__N_1412[28]), .CK(clk_N_875), .Q(multOut[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam multOut_i28.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_adj_70 (.A(n1068), .B(n3840), .C(n21440), .D(clk_N_875_enable_359), 
         .Z(n15130)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_70.init = 16'hfe00;
    LUT4 i3380_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m2[8]), .Z(n5882)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3380_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_adj_71 (.A(n16670), .B(n16296), .C(n21463), .D(n22216), 
         .Z(clk_N_875_enable_392)) /* synthesis lut_function=((B (C (D))+!B (C+!(D)))+!A) */ ;
    defparam i1_4_lut_adj_71.init = 16'hf577;
    LUT4 i1_2_lut_adj_72 (.A(Out2[8]), .B(Out2[12]), .Z(n6_adj_2339)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam i1_2_lut_adj_72.init = 16'heeee;
    LUT4 i1_4_lut_adj_73 (.A(n3704), .B(n35_adj_2340), .C(n40), .D(n36), 
         .Z(n4_adj_2341)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_73.init = 16'haaa8;
    LUT4 i14_4_lut (.A(speed_set_m3[13]), .B(speed_set_m3[1]), .C(speed_set_m3[12]), 
         .D(speed_set_m3[2]), .Z(n35_adj_2340)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(speed_set_m3[15]), .B(n38), .C(n32), .D(speed_set_m3[10]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i3384_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m2[10]), .Z(n5886)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3384_3_lut_4_lut.init = 16'hfd20;
    LUT4 i7_4_lut_adj_74 (.A(Out1[3]), .B(n14_adj_2342), .C(n10_adj_2343), 
         .D(Out1[4]), .Z(n18721)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i7_4_lut_adj_74.init = 16'hfffe;
    LUT4 i15_4_lut (.A(speed_set_m3[0]), .B(speed_set_m3[7]), .C(speed_set_m3[17]), 
         .D(speed_set_m3[11]), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(speed_set_m3[8]), .B(n34), .C(n24), .D(speed_set_m3[16]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut_adj_75 (.A(Out1[11]), .B(Out1[7]), .C(Out1[2]), .D(Out1[10]), 
         .Z(n14_adj_2342)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i6_4_lut_adj_75.init = 16'hfffe;
    LUT4 i11_3_lut (.A(speed_set_m3[6]), .B(speed_set_m3[3]), .C(speed_set_m3[14]), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut.init = 16'hfefe;
    LUT4 i2_2_lut_adj_76 (.A(Out1[9]), .B(Out1[1]), .Z(n10_adj_2343)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i2_2_lut_adj_76.init = 16'heeee;
    LUT4 i4_4_lut_adj_77 (.A(Out1[5]), .B(Out1[6]), .C(Out1[0]), .D(n6_adj_2344), 
         .Z(n18722)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i4_4_lut_adj_77.init = 16'hfffe;
    LUT4 i13_4_lut (.A(speed_set_m3[20]), .B(speed_set_m3[19]), .C(speed_set_m3[9]), 
         .D(speed_set_m3[4]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_78 (.A(Out1[8]), .B(Out1[12]), .Z(n6_adj_2344)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam i1_2_lut_adj_78.init = 16'heeee;
    LUT4 i3_2_lut_adj_79 (.A(speed_set_m3[18]), .B(speed_set_m3[5]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_79.init = 16'heeee;
    FD1P3AX Out0_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i1.GSR = "ENABLED";
    FD1P3AX Out0_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i2.GSR = "ENABLED";
    FD1P3AX Out0_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i3.GSR = "ENABLED";
    FD1P3AX Out0_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i4.GSR = "ENABLED";
    FD1P3AX Out0_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i5.GSR = "ENABLED";
    FD1P3AX Out0_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i6.GSR = "ENABLED";
    FD1P3AX Out0_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i7.GSR = "ENABLED";
    FD1P3AX Out0_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i8.GSR = "ENABLED";
    FD1P3AX Out0_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i9.GSR = "ENABLED";
    FD1P3AX Out0_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i10.GSR = "ENABLED";
    FD1P3AX Out0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i11.GSR = "ENABLED";
    FD1P3AX Out0_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i12.GSR = "ENABLED";
    FD1P3AX Out0_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i13.GSR = "ENABLED";
    FD1P3AX Out0_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i14.GSR = "ENABLED";
    FD1P3AX Out0_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i15.GSR = "ENABLED";
    FD1P3AX Out0_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i16.GSR = "ENABLED";
    FD1P3AX Out0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i17.GSR = "ENABLED";
    FD1P3AX Out0_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i18.GSR = "ENABLED";
    FD1P3AX Out0_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i19.GSR = "ENABLED";
    FD1P3AX Out0_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i20.GSR = "ENABLED";
    FD1P3AX Out0_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i21.GSR = "ENABLED";
    FD1P3AX Out0_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i22.GSR = "ENABLED";
    FD1P3AX Out0_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i23.GSR = "ENABLED";
    FD1P3AX Out0_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i24.GSR = "ENABLED";
    FD1P3AX Out0_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i25.GSR = "ENABLED";
    FD1P3AX Out0_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i26.GSR = "ENABLED";
    FD1P3AX Out0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i27.GSR = "ENABLED";
    FD1P3AX Out0_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_97), 
            .CK(clk_N_875), .Q(Out0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out0_i28.GSR = "ENABLED";
    FD1P3AX Out1_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i1.GSR = "ENABLED";
    FD1P3AX Out1_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i2.GSR = "ENABLED";
    FD1P3AX Out1_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i3.GSR = "ENABLED";
    FD1P3AX Out1_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i4.GSR = "ENABLED";
    FD1P3AX Out1_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i5.GSR = "ENABLED";
    FD1P3AX Out1_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i6.GSR = "ENABLED";
    FD1P3AX Out1_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i7.GSR = "ENABLED";
    FD1P3AX Out1_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i8.GSR = "ENABLED";
    FD1P3AX Out1_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i9.GSR = "ENABLED";
    FD1P3AX Out1_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i10.GSR = "ENABLED";
    FD1P3AX Out1_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i11.GSR = "ENABLED";
    FD1P3AX Out1_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i12.GSR = "ENABLED";
    FD1P3AX Out1_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i13.GSR = "ENABLED";
    FD1P3AX Out1_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i14.GSR = "ENABLED";
    FD1P3AX Out1_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i15.GSR = "ENABLED";
    FD1P3AX Out1_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i16.GSR = "ENABLED";
    FD1P3AX Out1_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i17.GSR = "ENABLED";
    FD1P3AX Out1_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i18.GSR = "ENABLED";
    FD1P3AX Out1_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i19.GSR = "ENABLED";
    FD1P3AX Out1_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i20.GSR = "ENABLED";
    FD1P3AX Out1_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i21.GSR = "ENABLED";
    FD1P3AX Out1_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i22.GSR = "ENABLED";
    FD1P3AX Out1_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i23.GSR = "ENABLED";
    FD1P3AX Out1_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i24.GSR = "ENABLED";
    FD1P3AX Out1_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i25.GSR = "ENABLED";
    FD1P3AX Out1_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i26.GSR = "ENABLED";
    FD1P3AX Out1_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i27.GSR = "ENABLED";
    FD1P3AX Out1_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_125), 
            .CK(clk_N_875), .Q(Out1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out1_i28.GSR = "ENABLED";
    FD1P3AX Out2_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i1.GSR = "ENABLED";
    FD1P3AX Out2_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i2.GSR = "ENABLED";
    FD1P3AX Out2_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i3.GSR = "ENABLED";
    FD1P3AX Out2_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i4.GSR = "ENABLED";
    FD1P3AX Out2_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i5.GSR = "ENABLED";
    FD1P3AX Out2_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i6.GSR = "ENABLED";
    FD1P3AX Out2_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i7.GSR = "ENABLED";
    FD1P3AX Out2_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i8.GSR = "ENABLED";
    FD1P3AX Out2_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i9.GSR = "ENABLED";
    FD1P3AX Out2_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i10.GSR = "ENABLED";
    FD1P3AX Out2_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i11.GSR = "ENABLED";
    FD1P3AX Out2_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i12.GSR = "ENABLED";
    FD1P3AX Out2_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i13.GSR = "ENABLED";
    FD1P3AX Out2_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i14.GSR = "ENABLED";
    FD1P3AX Out2_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i15.GSR = "ENABLED";
    FD1P3AX Out2_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i16.GSR = "ENABLED";
    FD1P3AX Out2_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i17.GSR = "ENABLED";
    FD1P3AX Out2_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i18.GSR = "ENABLED";
    FD1P3AX Out2_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i19.GSR = "ENABLED";
    FD1P3AX Out2_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i20.GSR = "ENABLED";
    FD1P3AX Out2_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i21.GSR = "ENABLED";
    FD1P3AX Out2_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i22.GSR = "ENABLED";
    FD1P3AX Out2_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i23.GSR = "ENABLED";
    FD1P3AX Out2_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i24.GSR = "ENABLED";
    FD1P3AX Out2_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i25.GSR = "ENABLED";
    FD1P3AX Out2_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i26.GSR = "ENABLED";
    FD1P3AX Out2_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i27.GSR = "ENABLED";
    FD1P3AX Out2_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_153), 
            .CK(clk_N_875), .Q(Out2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out2_i28.GSR = "ENABLED";
    FD1P3AX Out3_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i1.GSR = "ENABLED";
    FD1P3AX Out3_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i2.GSR = "ENABLED";
    FD1P3AX Out3_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i3.GSR = "ENABLED";
    FD1P3AX Out3_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i4.GSR = "ENABLED";
    FD1P3AX Out3_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i5.GSR = "ENABLED";
    FD1P3AX Out3_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i6.GSR = "ENABLED";
    FD1P3AX Out3_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i7.GSR = "ENABLED";
    FD1P3AX Out3_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i8.GSR = "ENABLED";
    FD1P3AX Out3_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i9.GSR = "ENABLED";
    FD1P3AX Out3_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i10.GSR = "ENABLED";
    FD1P3AX Out3_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i11.GSR = "ENABLED";
    FD1P3AX Out3_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i12.GSR = "ENABLED";
    FD1P3AX Out3_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i13.GSR = "ENABLED";
    FD1P3AX Out3_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i14.GSR = "ENABLED";
    FD1P3AX Out3_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i15.GSR = "ENABLED";
    FD1P3AX Out3_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i16.GSR = "ENABLED";
    FD1P3AX Out3_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i17.GSR = "ENABLED";
    FD1P3AX Out3_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i18.GSR = "ENABLED";
    FD1P3AX Out3_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i19.GSR = "ENABLED";
    FD1P3AX Out3_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i20.GSR = "ENABLED";
    FD1P3AX Out3_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i21.GSR = "ENABLED";
    FD1P3AX Out3_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i22.GSR = "ENABLED";
    FD1P3AX Out3_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i23.GSR = "ENABLED";
    FD1P3AX Out3_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i24.GSR = "ENABLED";
    FD1P3AX Out3_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i25.GSR = "ENABLED";
    FD1P3AX Out3_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i26.GSR = "ENABLED";
    FD1P3AX Out3_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i27.GSR = "ENABLED";
    FD1P3AX Out3_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_181), 
            .CK(clk_N_875), .Q(Out3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam Out3_i28.GSR = "ENABLED";
    FD1P3AX backOut2_i0_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut2_i0_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_209), 
            .CK(clk_N_875), .Q(backOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut2_i0_i28.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i1 (.D(backOut3_28__N_1874[1]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i1.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i2 (.D(backOut3_28__N_1874[2]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i2.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i3 (.D(backOut3_28__N_1874[3]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i3.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i4 (.D(backOut3_28__N_1874[4]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i4.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i5 (.D(backOut3_28__N_1874[5]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i5.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i6 (.D(backOut3_28__N_1874[6]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i6.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i7 (.D(backOut3_28__N_1874[7]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i7.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i8 (.D(backOut3_28__N_1874[8]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i8.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i9 (.D(backOut3_28__N_1874[9]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i9.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i10 (.D(backOut3_28__N_1874[10]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i10.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i11 (.D(Out2_28__N_1145[11]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i11.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i12 (.D(backOut3_28__N_1874[12]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i12.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i13 (.D(backOut3_28__N_1874[13]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i13.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i14 (.D(backOut3_28__N_1874[14]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i14.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i15 (.D(backOut3_28__N_1874[15]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i15.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i16 (.D(backOut3_28__N_1874[16]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i16.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i17 (.D(Out2_28__N_1145[17]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i17.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i18 (.D(backOut3_28__N_1874[18]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i18.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i19 (.D(Out2_28__N_1145[19]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i19.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i20 (.D(Out2_28__N_1145[20]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i20.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i21 (.D(backOut3_28__N_1874[21]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i21.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i22 (.D(backOut3_28__N_1874[22]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i22.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i23 (.D(backOut3_28__N_1874[23]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i23.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i24 (.D(Out2_28__N_1145[24]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i24.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i25 (.D(Out2_28__N_1145[25]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i25.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i26 (.D(Out0_28__N_1087[26]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i26.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i27 (.D(Out0_28__N_1087[27]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i27.GSR = "DISABLED";
    FD1P3AX backOut3_i0_i28 (.D(backOut2_28__N_1845[28]), .SP(clk_N_875_enable_237), 
            .CK(clk_N_875), .Q(backOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam backOut3_i0_i28.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_80 (.A(n16678), .B(n18698), .C(n21463), .D(n22216), 
         .Z(clk_N_875_enable_359)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;
    defparam i1_4_lut_adj_80.init = 16'hf5dd;
    LUT4 mux_92_i15_4_lut (.A(\speed_avg_m4[14] ), .B(\speed_avg_m3[14] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i15_4_lut.init = 16'hcac0;
    LUT4 mux_92_i14_4_lut (.A(\speed_avg_m4[13] ), .B(\speed_avg_m3[13] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i14_4_lut.init = 16'hcac0;
    LUT4 mux_92_i12_4_lut (.A(\speed_avg_m4[11] ), .B(\speed_avg_m3[11] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i12_4_lut.init = 16'hcac0;
    LUT4 mux_92_i11_4_lut (.A(\speed_avg_m4[10] ), .B(\speed_avg_m3[10] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i11_4_lut.init = 16'hcac0;
    FD1S3AX subOut_i1 (.D(\subOut_24__N_1369[1] ), .CK(clk_N_875), .Q(subOut[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i1.GSR = "ENABLED";
    FD1S3AX subOut_i2 (.D(\subOut_24__N_1369[2] ), .CK(clk_N_875), .Q(subOut[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i2.GSR = "ENABLED";
    FD1S3AX subOut_i3 (.D(\subOut_24__N_1369[3] ), .CK(clk_N_875), .Q(subOut[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i3.GSR = "ENABLED";
    FD1S3AX subOut_i4 (.D(\subOut_24__N_1369[4] ), .CK(clk_N_875), .Q(subOut[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i4.GSR = "ENABLED";
    FD1S3AX subOut_i5 (.D(\subOut_24__N_1369[5] ), .CK(clk_N_875), .Q(subOut[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i5.GSR = "ENABLED";
    FD1S3AX subOut_i6 (.D(\subOut_24__N_1369[6] ), .CK(clk_N_875), .Q(subOut[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i6.GSR = "ENABLED";
    FD1S3AX subOut_i7 (.D(\subOut_24__N_1369[7] ), .CK(clk_N_875), .Q(subOut[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i7.GSR = "ENABLED";
    FD1S3AX subOut_i8 (.D(\subOut_24__N_1369[8] ), .CK(clk_N_875), .Q(subOut[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i8.GSR = "ENABLED";
    FD1S3AX subOut_i9 (.D(\subOut_24__N_1369[9] ), .CK(clk_N_875), .Q(subOut[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i9.GSR = "ENABLED";
    FD1S3AX subOut_i10 (.D(\subOut_24__N_1369[10] ), .CK(clk_N_875), .Q(subOut[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i10.GSR = "ENABLED";
    FD1S3AX subOut_i11 (.D(\subOut_24__N_1369[11] ), .CK(clk_N_875), .Q(subOut[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i11.GSR = "ENABLED";
    FD1S3AX subOut_i12 (.D(\subOut_24__N_1369[12] ), .CK(clk_N_875), .Q(subOut[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i12.GSR = "ENABLED";
    FD1S3AX subOut_i13 (.D(\subOut_24__N_1369[13] ), .CK(clk_N_875), .Q(subOut[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i13.GSR = "ENABLED";
    FD1S3AX subOut_i14 (.D(\subOut_24__N_1369[14] ), .CK(clk_N_875), .Q(subOut[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i14.GSR = "ENABLED";
    FD1S3AX subOut_i15 (.D(\subOut_24__N_1369[15] ), .CK(clk_N_875), .Q(subOut[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i15.GSR = "ENABLED";
    FD1S3AX subOut_i16 (.D(\subOut_24__N_1369[16] ), .CK(clk_N_875), .Q(subOut[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i16.GSR = "ENABLED";
    FD1S3AX subOut_i17 (.D(\subOut_24__N_1369[17] ), .CK(clk_N_875), .Q(subOut[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i17.GSR = "ENABLED";
    FD1S3AX subOut_i18 (.D(\subOut_24__N_1369[18] ), .CK(clk_N_875), .Q(subOut[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i18.GSR = "ENABLED";
    FD1S3AX subOut_i19 (.D(\subOut_24__N_1369[19] ), .CK(clk_N_875), .Q(subOut[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i19.GSR = "ENABLED";
    FD1S3AX subOut_i20 (.D(\subOut_24__N_1369[20] ), .CK(clk_N_875), .Q(subOut[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i20.GSR = "ENABLED";
    FD1S3AX subOut_i21 (.D(\subOut_24__N_1369[21] ), .CK(clk_N_875), .Q(subOut[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i21.GSR = "ENABLED";
    FD1S3AX subOut_i23 (.D(\subOut_24__N_1369[24] ), .CK(clk_N_875), .Q(subOut[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam subOut_i23.GSR = "ENABLED";
    LUT4 mux_1221_i11_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[10]), 
         .D(speed_set_m4[10]), .Z(n5409)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_81 (.A(n3656), .B(n35_adj_2345), .C(n40_adj_2346), 
         .D(n36_adj_2347), .Z(n4_adj_2348)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_81.init = 16'haaa8;
    LUT4 mux_1221_i16_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m4[15]), .Z(n5419)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i14_4_lut_adj_82 (.A(speed_set_m2[13]), .B(speed_set_m2[1]), .C(speed_set_m2[12]), 
         .D(speed_set_m2[2]), .Z(n35_adj_2345)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_82.init = 16'hfffe;
    LUT4 mux_1221_i18_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m4[17]), .Z(n5423)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1221_i17_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m4[16]), .Z(n5421)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_92_i7_4_lut (.A(\speed_avg_m4[6] ), .B(\speed_avg_m3[6] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i7_4_lut.init = 16'hcac0;
    LUT4 mux_189_i22_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[21]), 
         .Z(intgOut0_28__N_1629[21])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i22_3_lut_3_lut.init = 16'hbaba;
    LUT4 i19_4_lut_adj_83 (.A(speed_set_m2[15]), .B(n38_adj_2349), .C(n32_adj_2350), 
         .D(speed_set_m2[10]), .Z(n40_adj_2346)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_83.init = 16'hfffe;
    LUT4 i15_4_lut_adj_84 (.A(speed_set_m2[0]), .B(speed_set_m2[7]), .C(speed_set_m2[17]), 
         .D(speed_set_m2[11]), .Z(n36_adj_2347)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_84.init = 16'hfffe;
    LUT4 i3386_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m2[11]), .Z(n5888)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3386_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i6_4_lut (.A(\speed_avg_m4[5] ), .B(\speed_avg_m3[5] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i6_4_lut.init = 16'hcac0;
    LUT4 i17_4_lut_adj_85 (.A(speed_set_m2[8]), .B(n34_adj_2351), .C(n24_adj_2352), 
         .D(speed_set_m2[16]), .Z(n38_adj_2349)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_85.init = 16'hfffe;
    LUT4 i11_3_lut_adj_86 (.A(speed_set_m2[6]), .B(speed_set_m2[3]), .C(speed_set_m2[14]), 
         .Z(n32_adj_2350)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_86.init = 16'hfefe;
    LUT4 mux_1221_i9_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[8]), 
         .D(speed_set_m4[8]), .Z(n5405)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_189_i20_3_lut_3_lut (.A(n1068), .B(n3840), .C(addOut[19]), 
         .Z(intgOut0_28__N_1629[19])) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam mux_189_i20_3_lut_3_lut.init = 16'hbaba;
    LUT4 mux_92_i5_4_lut (.A(\speed_avg_m4[4] ), .B(\speed_avg_m3[4] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i5_4_lut.init = 16'hcac0;
    LUT4 i13_4_lut_adj_87 (.A(speed_set_m2[20]), .B(speed_set_m2[19]), .C(speed_set_m2[9]), 
         .D(speed_set_m2[4]), .Z(n34_adj_2351)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_87.init = 16'hfffe;
    LUT4 i3_2_lut_adj_88 (.A(speed_set_m2[18]), .B(speed_set_m2[5]), .Z(n24_adj_2352)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_88.init = 16'heeee;
    LUT4 i3388_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[12]), 
         .D(speed_set_m2[12]), .Z(n5890)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3388_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_92_i3_4_lut (.A(\speed_avg_m4[2] ), .B(\speed_avg_m3[2] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i3_4_lut.init = 16'hcac0;
    LUT4 mux_92_i2_4_lut (.A(\speed_avg_m4[1] ), .B(\speed_avg_m3[1] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i2_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut_adj_89 (.A(n16301), .B(n19646), .C(n21463), .D(n22216), 
         .Z(clk_N_875_enable_387)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;
    defparam i1_4_lut_adj_89.init = 16'hf5dd;
    LUT4 mux_92_i1_4_lut (.A(\speed_avg_m4[0] ), .B(\speed_avg_m3[0] ), 
         .C(n21448), .D(n4389), .Z(subIn2_24__N_1535[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(147[18] 151[17])
    defparam mux_92_i1_4_lut.init = 16'hcac0;
    LUT4 mux_1221_i3_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[2]), 
         .D(speed_set_m4[2]), .Z(n5393)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_90 (.A(n16674), .B(n19672), .C(n21463), .D(n22216), 
         .Z(clk_N_875_enable_303)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;
    defparam i1_4_lut_adj_90.init = 16'hf5dd;
    LUT4 i1_4_lut_adj_91 (.A(n3608), .B(n35_adj_2353), .C(n40_adj_2354), 
         .D(n36_adj_2355), .Z(n4_adj_2356)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_91.init = 16'haaa8;
    LUT4 i14_4_lut_adj_92 (.A(speed_set_m1[13]), .B(speed_set_m1[1]), .C(speed_set_m1[12]), 
         .D(speed_set_m1[2]), .Z(n35_adj_2353)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i14_4_lut_adj_92.init = 16'hfffe;
    LUT4 i19_4_lut_adj_93 (.A(speed_set_m1[15]), .B(n38_adj_2357), .C(n32_adj_2358), 
         .D(speed_set_m1[10]), .Z(n40_adj_2354)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i19_4_lut_adj_93.init = 16'hfffe;
    LUT4 i15_4_lut_adj_94 (.A(speed_set_m1[0]), .B(speed_set_m1[7]), .C(speed_set_m1[17]), 
         .D(speed_set_m1[11]), .Z(n36_adj_2355)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i15_4_lut_adj_94.init = 16'hfffe;
    LUT4 mux_135_i22_4_lut (.A(backOut2[21]), .B(backOut3[21]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i22_4_lut.init = 16'h0aca;
    LUT4 i3390_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[13]), 
         .D(speed_set_m2[13]), .Z(n5892)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3390_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17_4_lut_adj_95 (.A(speed_set_m1[8]), .B(n34_adj_2359), .C(n24_adj_2360), 
         .D(speed_set_m1[16]), .Z(n38_adj_2357)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i17_4_lut_adj_95.init = 16'hfffe;
    LUT4 i1_4_lut_adj_96 (.A(n3752), .B(n35_adj_2361), .C(n40_adj_2362), 
         .D(n36_adj_2363), .Z(n4_adj_2364)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_96.init = 16'haaa8;
    LUT4 i14_4_lut_adj_97 (.A(speed_set_m4[13]), .B(speed_set_m4[1]), .C(speed_set_m4[12]), 
         .D(speed_set_m4[2]), .Z(n35_adj_2361)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut_adj_97.init = 16'hfffe;
    LUT4 i19_4_lut_adj_98 (.A(speed_set_m4[15]), .B(n38_adj_2365), .C(n32_adj_2366), 
         .D(speed_set_m4[10]), .Z(n40_adj_2362)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_98.init = 16'hfffe;
    LUT4 i15_4_lut_adj_99 (.A(speed_set_m4[0]), .B(speed_set_m4[7]), .C(speed_set_m4[17]), 
         .D(speed_set_m4[11]), .Z(n36_adj_2363)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_99.init = 16'hfffe;
    LUT4 i11_3_lut_adj_100 (.A(speed_set_m1[6]), .B(speed_set_m1[3]), .C(speed_set_m1[14]), 
         .Z(n32_adj_2358)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i11_3_lut_adj_100.init = 16'hfefe;
    LUT4 i17137_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21466), .D(n21467), .Z(n20157)) /* synthesis lut_function=(!((B (C (D))+!B (D))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(168[20:27])
    defparam i17137_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h08aa;
    LUT4 i17_4_lut_adj_101 (.A(speed_set_m4[8]), .B(n34_adj_2367), .C(n24_adj_2368), 
         .D(speed_set_m4[16]), .Z(n38_adj_2365)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_101.init = 16'hfffe;
    LUT4 i3392_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m2[14]), .Z(n5894)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3392_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13_4_lut_adj_102 (.A(speed_set_m1[20]), .B(speed_set_m1[19]), 
         .C(speed_set_m1[9]), .D(speed_set_m1[4]), .Z(n34_adj_2359)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i13_4_lut_adj_102.init = 16'hfffe;
    LUT4 i11_3_lut_adj_103 (.A(speed_set_m4[6]), .B(speed_set_m4[3]), .C(speed_set_m4[14]), 
         .Z(n32_adj_2366)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11_3_lut_adj_103.init = 16'hfefe;
    LUT4 i13_4_lut_adj_104 (.A(speed_set_m4[20]), .B(speed_set_m4[19]), 
         .C(speed_set_m4[9]), .D(speed_set_m4[4]), .Z(n34_adj_2367)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_104.init = 16'hfffe;
    LUT4 i3_2_lut_adj_105 (.A(speed_set_m4[18]), .B(speed_set_m4[5]), .Z(n24_adj_2368)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_adj_105.init = 16'heeee;
    LUT4 mux_135_i23_4_lut (.A(backOut2[22]), .B(backOut3[22]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i23_4_lut.init = 16'h0aca;
    LUT4 mux_135_i2_4_lut (.A(backOut2[1]), .B(backOut3[1]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i2_4_lut.init = 16'h0aca;
    LUT4 mux_135_i24_4_lut (.A(backOut2[23]), .B(backOut3[23]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i24_4_lut.init = 16'h0aca;
    LUT4 mux_135_i3_4_lut (.A(backOut2[2]), .B(backOut3[2]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i3_4_lut.init = 16'h0aca;
    LUT4 mux_135_i25_4_lut (.A(backOut2[24]), .B(backOut3[24]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i25_4_lut.init = 16'h0aca;
    LUT4 mux_135_i4_4_lut (.A(backOut2[3]), .B(backOut3[3]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i4_4_lut.init = 16'h0aca;
    LUT4 mux_135_i26_4_lut (.A(backOut2[25]), .B(backOut3[25]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i26_4_lut.init = 16'h0aca;
    LUT4 mux_135_i5_4_lut (.A(backOut2[4]), .B(backOut3[4]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i5_4_lut.init = 16'h0aca;
    LUT4 mux_135_i27_4_lut (.A(backOut2[26]), .B(backOut3[26]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i27_4_lut.init = 16'h0aca;
    LUT4 mux_135_i6_4_lut (.A(backOut2[5]), .B(backOut3[5]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i6_4_lut.init = 16'h0aca;
    LUT4 i17235_2_lut_3_lut_4_lut (.A(n21430), .B(n21418), .C(multIn2[11]), 
         .D(multIn2[0]), .Z(multIn2[9])) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam i17235_2_lut_3_lut_4_lut.init = 16'hf0f7;
    LUT4 mux_135_i7_4_lut (.A(backOut2[6]), .B(backOut3[6]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i7_4_lut.init = 16'h0aca;
    LUT4 mux_135_i28_4_lut (.A(backOut2[27]), .B(backOut3[27]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i28_4_lut.init = 16'h0aca;
    LUT4 mux_135_i8_4_lut (.A(backOut2[7]), .B(backOut3[7]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i8_4_lut.init = 16'h0aca;
    LUT4 i7_4_lut_adj_106 (.A(Out0[3]), .B(n14_adj_2369), .C(n10_adj_2370), 
         .D(Out0[4]), .Z(n18759)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i7_4_lut_adj_106.init = 16'hfffe;
    LUT4 i6_4_lut_adj_107 (.A(Out0[11]), .B(Out0[7]), .C(Out0[2]), .D(Out0[10]), 
         .Z(n14_adj_2369)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i6_4_lut_adj_107.init = 16'hfffe;
    LUT4 i2_2_lut_adj_108 (.A(Out0[9]), .B(Out0[1]), .Z(n10_adj_2370)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i2_2_lut_adj_108.init = 16'heeee;
    LUT4 i4_4_lut_adj_109 (.A(Out0[5]), .B(Out0[6]), .C(Out0[0]), .D(n6_adj_2371), 
         .Z(n18760)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i4_4_lut_adj_109.init = 16'hfffe;
    LUT4 i1_2_lut_adj_110 (.A(Out0[8]), .B(Out0[12]), .Z(n6_adj_2371)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam i1_2_lut_adj_110.init = 16'heeee;
    LUT4 mux_135_i29_4_lut (.A(backOut2[28]), .B(backOut3[28]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i29_4_lut.init = 16'h0aca;
    LUT4 mux_135_i9_4_lut (.A(backOut2[8]), .B(backOut3[8]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i9_4_lut.init = 16'h0aca;
    LUT4 mux_135_i10_4_lut (.A(backOut2[9]), .B(backOut3[9]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i10_4_lut.init = 16'h0aca;
    LUT4 mux_135_i11_4_lut (.A(backOut2[10]), .B(backOut3[10]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i11_4_lut.init = 16'h0aca;
    LUT4 mux_135_i12_4_lut (.A(backOut2[11]), .B(backOut3[11]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i12_4_lut.init = 16'h0aca;
    LUT4 mux_135_i13_4_lut (.A(backOut2[12]), .B(backOut3[12]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i13_4_lut.init = 16'h0aca;
    LUT4 mux_135_i14_4_lut (.A(backOut2[13]), .B(backOut3[13]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i14_4_lut.init = 16'h0aca;
    LUT4 mux_135_i15_4_lut (.A(backOut2[14]), .B(backOut3[14]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i15_4_lut.init = 16'h0aca;
    LUT4 mux_135_i16_4_lut (.A(backOut2[15]), .B(backOut3[15]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i16_4_lut.init = 16'h0aca;
    LUT4 mux_135_i17_4_lut (.A(backOut2[16]), .B(backOut3[16]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i17_4_lut.init = 16'h0aca;
    LUT4 mux_1221_i12_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[11]), 
         .D(speed_set_m4[11]), .Z(n5411)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_135_i18_4_lut (.A(backOut2[17]), .B(backOut3[17]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i18_4_lut.init = 16'h0aca;
    LUT4 i3_2_lut_adj_111 (.A(speed_set_m1[18]), .B(speed_set_m1[5]), .Z(n24_adj_2360)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[7:22])
    defparam i3_2_lut_adj_111.init = 16'heeee;
    LUT4 mux_91_i13_3_lut_4_lut_4_lut (.A(n21420), .B(\speed_avg_m4[12] ), 
         .C(n4389), .D(n21418), .Z(n367[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i13_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_135_i19_4_lut (.A(backOut2[18]), .B(backOut3[18]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i19_4_lut.init = 16'h0aca;
    LUT4 mux_91_i10_3_lut_4_lut_4_lut (.A(n21420), .B(\speed_avg_m4[9] ), 
         .C(n4389), .D(n21418), .Z(n367[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i10_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_135_i20_4_lut (.A(backOut2[19]), .B(backOut3[19]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i20_4_lut.init = 16'h0aca;
    LUT4 mux_91_i9_3_lut_4_lut_4_lut (.A(n21420), .B(\speed_avg_m4[8] ), 
         .C(n4389), .D(n21418), .Z(n367[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i9_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_91_i8_3_lut_4_lut_4_lut (.A(n21420), .B(\speed_avg_m4[7] ), 
         .C(n4389), .D(n21418), .Z(n367[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i8_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_91_i4_3_lut_4_lut_4_lut (.A(n21420), .B(\speed_avg_m4[3] ), 
         .C(n4389), .D(n21418), .Z(n367[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(171[9:16])
    defparam mux_91_i4_3_lut_4_lut_4_lut.init = 16'hcacf;
    LUT4 mux_135_i21_4_lut (.A(backOut2[20]), .B(backOut3[20]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i21_4_lut.init = 16'h0aca;
    LUT4 mux_135_i1_4_lut (.A(backOut2[0]), .B(backOut3[0]), .C(n21430), 
         .D(n9_adj_2327), .Z(n558[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 191[27])
    defparam mux_135_i1_4_lut.init = 16'h0aca;
    LUT4 i3394_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[15]), 
         .D(speed_set_m2[15]), .Z(n5896)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3394_3_lut_4_lut.init = 16'hfd20;
    LUT4 i17143_4_lut_4_lut (.A(n21446), .B(n20118), .C(n21444), .D(n21432), 
         .Z(n20127)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(184[17] 185[26])
    defparam i17143_4_lut_4_lut.init = 16'hdfff;
    LUT4 i1755_1_lut (.A(n42), .Z(subIn1_24__N_1534)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(137[34:50])
    defparam i1755_1_lut.init = 16'h5555;
    LUT4 i3396_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[16]), 
         .D(speed_set_m2[16]), .Z(n5898)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3396_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3398_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[17]), 
         .D(speed_set_m2[17]), .Z(n5900)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3398_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_323_3_lut_4_lut (.A(ss[2]), .B(n21475), .C(ss[1]), 
         .D(n22216), .Z(n21424)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_323_3_lut_4_lut.init = 16'hffef;
    LUT4 i3400_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m2[18]), .Z(n5902)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3400_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_326_3_lut_4_lut (.A(ss[2]), .B(n21475), .C(ss[1]), 
         .D(n22216), .Z(n21427)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_326_3_lut_4_lut.init = 16'hfffe;
    LUT4 i11718_2_lut_3_lut_4_lut (.A(n21494), .B(n21491), .C(clk_N_875_enable_387), 
         .D(ss[1]), .Z(n14304)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i11718_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i11746_2_lut_3_lut_4_lut (.A(n21494), .B(n21491), .C(clk_N_875_enable_359), 
         .D(ss[1]), .Z(n14332)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i11746_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i3402_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m2[19]), .Z(n5904)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3402_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2_3_lut_4_lut_adj_112 (.A(ss[1]), .B(n21493), .C(n22216), .D(ss[3]), 
         .Z(n19674)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_3_lut_4_lut_adj_112.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_113 (.A(n21492), .B(n21491), .C(n22211), 
         .D(n22216), .Z(n19662)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_113.init = 16'he0f0;
    LUT4 i1756_1_lut (.A(n49), .Z(dirout_m3_N_1949)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(139[35:51])
    defparam i1756_1_lut.init = 16'h5555;
    LUT4 i1754_1_lut (.A(n35), .Z(subIn1_24__N_1347)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(135[34:50])
    defparam i1754_1_lut.init = 16'h5555;
    LUT4 i1757_1_lut (.A(n56), .Z(dirout_m4_N_1952)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(141[35:51])
    defparam i1757_1_lut.init = 16'h5555;
    LUT4 i13373_2_lut (.A(addOut[28]), .B(n22216), .Z(backOut2_28__N_1845[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13373_2_lut.init = 16'h2222;
    LUT4 i13533_2_lut (.A(addOut[27]), .B(n22216), .Z(Out0_28__N_1087[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13533_2_lut.init = 16'h2222;
    LUT4 i13526_2_lut (.A(addOut[26]), .B(n22216), .Z(Out0_28__N_1087[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13526_2_lut.init = 16'h2222;
    LUT4 i13622_2_lut (.A(addOut[25]), .B(n22216), .Z(Out2_28__N_1145[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13622_2_lut.init = 16'h2222;
    LUT4 n15710_bdd_4_lut_rep_400 (.A(n21499), .B(ss[0]), .C(n22209), 
         .D(ss[1]), .Z(n22204)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam n15710_bdd_4_lut_rep_400.init = 16'h0410;
    LUT4 i17231_2_lut_3_lut_4_lut (.A(n21499), .B(n22203), .C(n22204), 
         .D(ss[2]), .Z(n20388)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i17231_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i3406_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m2[20]), .Z(n5908)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i3406_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_371 (.A(ss[1]), .B(ss[2]), .Z(n21472)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_371.init = 16'h2222;
    LUT4 i13150_2_lut_rep_372 (.A(ss[0]), .B(ss[1]), .Z(n21473)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13150_2_lut_rep_372.init = 16'h8888;
    LUT4 mux_1221_i2_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[1]), 
         .D(speed_set_m4[1]), .Z(n5391)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i7984_2_lut_3_lut (.A(ss[0]), .B(ss[1]), .C(ss[2]), .Z(n14)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i7984_2_lut_3_lut.init = 16'h7878;
    LUT4 ss_4__I_0_357_i9_2_lut_rep_345_3_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21498), .D(ss[3]), .Z(n21446)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam ss_4__I_0_357_i9_2_lut_rep_345_3_lut_4_lut.init = 16'hfff7;
    LUT4 ss_4__I_0_360_i9_2_lut_rep_343_3_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21494), .D(ss[3]), .Z(n21444)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam ss_4__I_0_360_i9_2_lut_rep_343_3_lut_4_lut.init = 16'hfff7;
    LUT4 equal_110_i9_2_lut_rep_342_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(n21498), 
         .D(ss[3]), .Z(n21443)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam equal_110_i9_2_lut_rep_342_3_lut_4_lut.init = 16'hf7ff;
    LUT4 mux_1221_i1_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[0]), 
         .D(speed_set_m4[0]), .Z(n5347)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_373 (.A(ss[2]), .B(ss[1]), .Z(n21474)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_373.init = 16'h2222;
    CCU2D add_1212_5 (.A0(n5439), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5441), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18232), 
          .COUT(n18233), .S0(n2373[3]), .S1(n2373[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_5.INIT0 = 16'hf555;
    defparam add_1212_5.INIT1 = 16'hf555;
    defparam add_1212_5.INJECT1_0 = "NO";
    defparam add_1212_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_374 (.A(ss[0]), .B(ss[3]), .Z(n21475)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_374.init = 16'hbbbb;
    LUT4 i2_2_lut_rep_357_3_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n21458)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i2_2_lut_rep_357_3_lut.init = 16'hfbfb;
    CCU2D add_223_13 (.A0(Out3[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18271), 
          .COUT(n18272), .S0(n1364[11]), .S1(n1364[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_13.INIT0 = 16'h5aaa;
    defparam add_223_13.INIT1 = 16'h5aaa;
    defparam add_223_13.INJECT1_0 = "NO";
    defparam add_223_13.INJECT1_1 = "NO";
    CCU2D add_223_11 (.A0(Out3[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18270), 
          .COUT(n18271), .S0(n1364[9]), .S1(n1364[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_11.INIT0 = 16'h5aaa;
    defparam add_223_11.INIT1 = 16'h5aaa;
    defparam add_223_11.INJECT1_0 = "NO";
    defparam add_223_11.INJECT1_1 = "NO";
    CCU2D add_1212_3 (.A0(n5435), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5437), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18231), 
          .COUT(n18232), .S0(n2373[1]), .S1(n2373[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_3.INIT0 = 16'hf555;
    defparam add_1212_3.INIT1 = 16'hf555;
    defparam add_1212_3.INJECT1_0 = "NO";
    defparam add_1212_3.INJECT1_1 = "NO";
    LUT4 mux_1221_i6_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[5]), 
         .D(speed_set_m4[5]), .Z(n5399)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i6_3_lut_4_lut.init = 16'hf780;
    CCU2D add_15127_25 (.A0(addOut[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18459), .COUT(n18460));
    defparam add_15127_25.INIT0 = 16'h0aaa;
    defparam add_15127_25.INIT1 = 16'h0aaa;
    defparam add_15127_25.INJECT1_0 = "NO";
    defparam add_15127_25.INJECT1_1 = "NO";
    CCU2D add_15127_23 (.A0(addOut[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18458), .COUT(n18459));
    defparam add_15127_23.INIT0 = 16'h0aaa;
    defparam add_15127_23.INIT1 = 16'h0aaa;
    defparam add_15127_23.INJECT1_0 = "NO";
    defparam add_15127_23.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut (.A(ss[0]), .B(ss[3]), .C(ss[2]), .Z(n19679)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut.init = 16'hbfbf;
    CCU2D add_1209_7 (.A0(n1364[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1364[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18336), 
          .COUT(n18337), .S0(n2317[5]), .S1(n2317[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1209_7.INIT0 = 16'hf555;
    defparam add_1209_7.INIT1 = 16'hf555;
    defparam add_1209_7.INJECT1_0 = "NO";
    defparam add_1209_7.INJECT1_1 = "NO";
    LUT4 i13711_2_lut_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), .D(n22209), 
         .Z(n16296)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13711_2_lut_3_lut_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_114 (.A(ss[0]), .B(ss[3]), .C(n22209), 
         .D(ss[1]), .Z(n19672)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_3_lut_4_lut_adj_114.init = 16'h0400;
    CCU2D add_1209_5 (.A0(n1364[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1364[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18335), 
          .COUT(n18336), .S0(n2317[3]), .S1(n2317[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1209_5.INIT0 = 16'hf555;
    defparam add_1209_5.INIT1 = 16'hf555;
    defparam add_1209_5.INJECT1_0 = "NO";
    defparam add_1209_5.INJECT1_1 = "NO";
    CCU2D add_15127_21 (.A0(addOut[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18457), .COUT(n18458));
    defparam add_15127_21.INIT0 = 16'h0aaa;
    defparam add_15127_21.INIT1 = 16'hf555;
    defparam add_15127_21.INJECT1_0 = "NO";
    defparam add_15127_21.INJECT1_1 = "NO";
    LUT4 i13617_2_lut (.A(addOut[24]), .B(n22216), .Z(Out2_28__N_1145[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13617_2_lut.init = 16'h2222;
    CCU2D add_15127_19 (.A0(addOut[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18456), .COUT(n18457));
    defparam add_15127_19.INIT0 = 16'hf555;
    defparam add_15127_19.INIT1 = 16'hf555;
    defparam add_15127_19.INJECT1_0 = "NO";
    defparam add_15127_19.INJECT1_1 = "NO";
    CCU2D add_1212_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5433), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18231), 
          .S1(n2373[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_1.INIT0 = 16'hF000;
    defparam add_1212_1.INIT1 = 16'h0aaa;
    defparam add_1212_1.INJECT1_0 = "NO";
    defparam add_1212_1.INJECT1_1 = "NO";
    LUT4 i2984_2_lut_rep_377 (.A(n22216), .B(n22211), .Z(clk_N_875_enable_391)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i2984_2_lut_rep_377.init = 16'h8888;
    LUT4 i11838_2_lut_3_lut_4_lut (.A(n22216), .B(n22211), .C(n21491), 
         .D(n21492), .Z(n14414)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11838_2_lut_3_lut_4_lut.init = 16'h8880;
    CCU2D add_15127_17 (.A0(addOut[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18455), .COUT(n18456));
    defparam add_15127_17.INIT0 = 16'hf555;
    defparam add_15127_17.INIT1 = 16'h0aaa;
    defparam add_15127_17.INJECT1_0 = "NO";
    defparam add_15127_17.INJECT1_1 = "NO";
    CCU2D add_1209_3 (.A0(n1364[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1364[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18334), 
          .COUT(n18335), .S0(n2317[1]), .S1(n2317[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1209_3.INIT0 = 16'hf555;
    defparam add_1209_3.INIT1 = 16'hf555;
    defparam add_1209_3.INJECT1_0 = "NO";
    defparam add_1209_3.INJECT1_1 = "NO";
    CCU2D add_15127_15 (.A0(addOut[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18454), .COUT(n18455));
    defparam add_15127_15.INIT0 = 16'hf555;
    defparam add_15127_15.INIT1 = 16'hf555;
    defparam add_15127_15.INJECT1_0 = "NO";
    defparam add_15127_15.INJECT1_1 = "NO";
    LUT4 i13728_2_lut_rep_305 (.A(n15757), .B(n56), .Z(n21406)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13728_2_lut_rep_305.init = 16'heeee;
    LUT4 mux_1222_i12_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[11]), 
         .D(speed_set_m3[11]), .Z(n5369)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3_2_lut_3_lut (.A(n15757), .B(n56), .C(subIn1_24__N_1342), .Z(n8_adj_2372)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;
    defparam i3_2_lut_3_lut.init = 16'h0e0e;
    LUT4 i14068_3_lut_4_lut (.A(n21465), .B(n21466), .C(n4_adj_2348), 
         .D(n3680), .Z(n16678)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i14068_3_lut_4_lut.init = 16'hfeee;
    LUT4 i13436_2_lut (.A(addOut[23]), .B(n22216), .Z(backOut3_28__N_1874[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13436_2_lut.init = 16'h2222;
    LUT4 i13433_2_lut (.A(addOut[22]), .B(n22216), .Z(backOut3_28__N_1874[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13433_2_lut.init = 16'h2222;
    LUT4 i13432_2_lut (.A(addOut[21]), .B(n22216), .Z(backOut3_28__N_1874[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13432_2_lut.init = 16'h2222;
    LUT4 i13610_2_lut (.A(addOut[20]), .B(n22216), .Z(Out2_28__N_1145[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13610_2_lut.init = 16'h2222;
    LUT4 i13609_2_lut (.A(addOut[19]), .B(n22216), .Z(Out2_28__N_1145[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13609_2_lut.init = 16'h2222;
    LUT4 i17264_2_lut_3_lut_3_lut_4_lut (.A(n21465), .B(n21464), .C(n21418), 
         .D(n21431), .Z(multIn2[3])) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(175[9:17])
    defparam i17264_2_lut_3_lut_3_lut_4_lut.init = 16'h001f;
    LUT4 i13419_2_lut (.A(addOut[18]), .B(n22216), .Z(backOut3_28__N_1874[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13419_2_lut.init = 16'h2222;
    CCU2D add_15127_13 (.A0(addOut[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18453), .COUT(n18454));
    defparam add_15127_13.INIT0 = 16'h0aaa;
    defparam add_15127_13.INIT1 = 16'h0aaa;
    defparam add_15127_13.INJECT1_0 = "NO";
    defparam add_15127_13.INJECT1_1 = "NO";
    CCU2D add_15127_11 (.A0(addOut[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18452), .COUT(n18453));
    defparam add_15127_11.INIT0 = 16'hf555;
    defparam add_15127_11.INIT1 = 16'h0aaa;
    defparam add_15127_11.INJECT1_0 = "NO";
    defparam add_15127_11.INJECT1_1 = "NO";
    CCU2D add_15127_9 (.A0(addOut[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18451), .COUT(n18452));
    defparam add_15127_9.INIT0 = 16'h0aaa;
    defparam add_15127_9.INIT1 = 16'hf555;
    defparam add_15127_9.INJECT1_0 = "NO";
    defparam add_15127_9.INJECT1_1 = "NO";
    CCU2D add_15127_7 (.A0(addOut[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18450), .COUT(n18451));
    defparam add_15127_7.INIT0 = 16'h0aaa;
    defparam add_15127_7.INIT1 = 16'hf555;
    defparam add_15127_7.INJECT1_0 = "NO";
    defparam add_15127_7.INJECT1_1 = "NO";
    CCU2D add_15127_5 (.A0(addOut[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18449), .COUT(n18450));
    defparam add_15127_5.INIT0 = 16'hf555;
    defparam add_15127_5.INIT1 = 16'hf555;
    defparam add_15127_5.INJECT1_0 = "NO";
    defparam add_15127_5.INJECT1_1 = "NO";
    CCU2D add_15127_3 (.A0(addOut[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18448), .COUT(n18449));
    defparam add_15127_3.INIT0 = 16'hf555;
    defparam add_15127_3.INIT1 = 16'hf555;
    defparam add_15127_3.INJECT1_0 = "NO";
    defparam add_15127_3.INJECT1_1 = "NO";
    CCU2D add_15127_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(addOut[0]), .B1(addOut[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18448));
    defparam add_15127_1.INIT0 = 16'hF000;
    defparam add_15127_1.INIT1 = 16'ha666;
    defparam add_15127_1.INJECT1_0 = "NO";
    defparam add_15127_1.INJECT1_1 = "NO";
    CCU2D add_15135_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18447), 
          .S0(n3632));
    defparam add_15135_cout.INIT0 = 16'h0000;
    defparam add_15135_cout.INIT1 = 16'h0000;
    defparam add_15135_cout.INJECT1_0 = "NO";
    defparam add_15135_cout.INJECT1_1 = "NO";
    CCU2D add_1209_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1364[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18334), 
          .S1(n2317[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(371[20:29])
    defparam add_1209_1.INIT0 = 16'hF000;
    defparam add_1209_1.INIT1 = 16'h0aaa;
    defparam add_1209_1.INJECT1_0 = "NO";
    defparam add_1209_1.INJECT1_1 = "NO";
    CCU2D add_15135_20 (.A0(speed_set_m1[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18446), .COUT(n18447));
    defparam add_15135_20.INIT0 = 16'h5aaa;
    defparam add_15135_20.INIT1 = 16'h0aaa;
    defparam add_15135_20.INJECT1_0 = "NO";
    defparam add_15135_20.INJECT1_1 = "NO";
    CCU2D add_15135_18 (.A0(speed_set_m1[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18445), .COUT(n18446));
    defparam add_15135_18.INIT0 = 16'h5aaa;
    defparam add_15135_18.INIT1 = 16'h5aaa;
    defparam add_15135_18.INJECT1_0 = "NO";
    defparam add_15135_18.INJECT1_1 = "NO";
    CCU2D add_1206_11 (.A0(n1301[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18230), 
          .S0(n2281[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1206_11.INIT0 = 16'hf555;
    defparam add_1206_11.INIT1 = 16'h0000;
    defparam add_1206_11.INJECT1_0 = "NO";
    defparam add_1206_11.INJECT1_1 = "NO";
    CCU2D add_1206_9 (.A0(n1301[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1301[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18229), 
          .COUT(n18230), .S0(n2281[7]), .S1(n2281[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1206_9.INIT0 = 16'hf555;
    defparam add_1206_9.INIT1 = 16'hf555;
    defparam add_1206_9.INJECT1_0 = "NO";
    defparam add_1206_9.INJECT1_1 = "NO";
    LUT4 i13726_2_lut_rep_306 (.A(n15773), .B(n49), .Z(n21407)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13726_2_lut_rep_306.init = 16'heeee;
    LUT4 i13607_2_lut (.A(addOut[17]), .B(n22216), .Z(Out2_28__N_1145[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13607_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_adj_115 (.A(n1343[15]), .B(n2305[8]), .C(n9_adj_2373), 
         .Z(n1502[8])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_115.init = 16'h8a8a;
    LUT4 mux_138_i2_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[1]), 
         .D(intgOut2[1]), .Z(n648[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i2_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1208_11 (.A0(n1343[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18333), 
          .S0(n2305[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1208_11.INIT0 = 16'hf555;
    defparam add_1208_11.INIT1 = 16'h0000;
    defparam add_1208_11.INJECT1_0 = "NO";
    defparam add_1208_11.INJECT1_1 = "NO";
    LUT4 mux_138_i22_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[21]), 
         .D(intgOut2[21]), .Z(n648[21])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i22_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i16_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[15]), 
         .D(intgOut2[15]), .Z(n648[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i16_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i11_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[10]), 
         .D(intgOut2[10]), .Z(n648[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i11_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_223_9 (.A0(Out3[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18269), 
          .COUT(n18270), .S0(n1364[7]), .S1(n1364[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_9.INIT0 = 16'h5aaa;
    defparam add_223_9.INIT1 = 16'h5aaa;
    defparam add_223_9.INJECT1_0 = "NO";
    defparam add_223_9.INJECT1_1 = "NO";
    LUT4 mux_138_i27_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[26]), 
         .D(intgOut2[26]), .Z(n648[26])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i27_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_rep_304_3_lut_4_lut (.A(n15773), .B(n49), .C(n56), .D(n15757), 
         .Z(n21405)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i1_2_lut_rep_304_3_lut_4_lut.init = 16'heee0;
    CCU2D add_223_7 (.A0(Out3[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18268), 
          .COUT(n18269), .S0(n1364[5]), .S1(n1364[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_7.INIT0 = 16'h5aaa;
    defparam add_223_7.INIT1 = 16'h5aaa;
    defparam add_223_7.INJECT1_0 = "NO";
    defparam add_223_7.INJECT1_1 = "NO";
    CCU2D add_223_5 (.A0(Out3[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18267), 
          .COUT(n18268), .S0(n1364[3]), .S1(n1364[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_5.INIT0 = 16'h5aaa;
    defparam add_223_5.INIT1 = 16'h5aaa;
    defparam add_223_5.INJECT1_0 = "NO";
    defparam add_223_5.INJECT1_1 = "NO";
    LUT4 mux_138_i26_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[25]), 
         .D(intgOut2[25]), .Z(n648[25])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i26_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1206_7 (.A0(n1301[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1301[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18228), 
          .COUT(n18229), .S0(n2281[5]), .S1(n2281[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1206_7.INIT0 = 16'hf555;
    defparam add_1206_7.INIT1 = 16'hf555;
    defparam add_1206_7.INJECT1_0 = "NO";
    defparam add_1206_7.INJECT1_1 = "NO";
    CCU2D add_223_3 (.A0(Out3[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18266), 
          .COUT(n18267), .S0(n1364[1]), .S1(n1364[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_3.INIT0 = 16'h5aaa;
    defparam add_223_3.INIT1 = 16'h5aaa;
    defparam add_223_3.INJECT1_0 = "NO";
    defparam add_223_3.INJECT1_1 = "NO";
    CCU2D add_1208_9 (.A0(n1343[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1343[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18332), 
          .COUT(n18333), .S0(n2305[7]), .S1(n2305[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1208_9.INIT0 = 16'hf555;
    defparam add_1208_9.INIT1 = 16'hf555;
    defparam add_1208_9.INJECT1_0 = "NO";
    defparam add_1208_9.INJECT1_1 = "NO";
    CCU2D add_1208_7 (.A0(n1343[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1343[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18331), 
          .COUT(n18332), .S0(n2305[5]), .S1(n2305[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1208_7.INIT0 = 16'hf555;
    defparam add_1208_7.INIT1 = 16'hf555;
    defparam add_1208_7.INJECT1_0 = "NO";
    defparam add_1208_7.INJECT1_1 = "NO";
    CCU2D add_1208_5 (.A0(n1343[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1343[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18330), 
          .COUT(n18331), .S0(n2305[3]), .S1(n2305[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1208_5.INIT0 = 16'hf555;
    defparam add_1208_5.INIT1 = 16'hf555;
    defparam add_1208_5.INJECT1_0 = "NO";
    defparam add_1208_5.INJECT1_1 = "NO";
    CCU2D add_1208_3 (.A0(n1343[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1343[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18329), 
          .COUT(n18330), .S0(n2305[1]), .S1(n2305[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1208_3.INIT0 = 16'hf555;
    defparam add_1208_3.INIT1 = 16'hf555;
    defparam add_1208_3.INJECT1_0 = "NO";
    defparam add_1208_3.INJECT1_1 = "NO";
    CCU2D add_15135_16 (.A0(speed_set_m1[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18444), .COUT(n18445));
    defparam add_15135_16.INIT0 = 16'h5aaa;
    defparam add_15135_16.INIT1 = 16'h5aaa;
    defparam add_15135_16.INJECT1_0 = "NO";
    defparam add_15135_16.INJECT1_1 = "NO";
    CCU2D add_223_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out3[13]), .B1(n18754), .C1(n18755), .D1(Out3[28]), .COUT(n18266), 
          .S1(n1364[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(337[17:21])
    defparam add_223_1.INIT0 = 16'hF000;
    defparam add_223_1.INIT1 = 16'h56aa;
    defparam add_223_1.INJECT1_0 = "NO";
    defparam add_223_1.INJECT1_1 = "NO";
    CCU2D add_219_17 (.A0(Out2[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18265), 
          .S0(n1343[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_17.INIT0 = 16'h5aaa;
    defparam add_219_17.INIT1 = 16'h0000;
    defparam add_219_17.INJECT1_0 = "NO";
    defparam add_219_17.INJECT1_1 = "NO";
    CCU2D add_219_15 (.A0(Out2[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18264), 
          .COUT(n18265), .S0(n1343[13]), .S1(n1343[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_15.INIT0 = 16'h5aaa;
    defparam add_219_15.INIT1 = 16'h5aaa;
    defparam add_219_15.INJECT1_0 = "NO";
    defparam add_219_15.INJECT1_1 = "NO";
    CCU2D add_219_13 (.A0(Out2[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18263), 
          .COUT(n18264), .S0(n1343[11]), .S1(n1343[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_13.INIT0 = 16'h5aaa;
    defparam add_219_13.INIT1 = 16'h5aaa;
    defparam add_219_13.INJECT1_0 = "NO";
    defparam add_219_13.INJECT1_1 = "NO";
    CCU2D add_219_11 (.A0(Out2[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18262), 
          .COUT(n18263), .S0(n1343[9]), .S1(n1343[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_11.INIT0 = 16'h5aaa;
    defparam add_219_11.INIT1 = 16'h5aaa;
    defparam add_219_11.INJECT1_0 = "NO";
    defparam add_219_11.INJECT1_1 = "NO";
    CCU2D add_1208_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1343[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18329), 
          .S1(n2305[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(363[20:29])
    defparam add_1208_1.INIT0 = 16'hF000;
    defparam add_1208_1.INIT1 = 16'h0aaa;
    defparam add_1208_1.INJECT1_0 = "NO";
    defparam add_1208_1.INJECT1_1 = "NO";
    CCU2D add_1207_11 (.A0(n1322[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18328), 
          .S0(n2293[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1207_11.INIT0 = 16'hf555;
    defparam add_1207_11.INIT1 = 16'h0000;
    defparam add_1207_11.INJECT1_0 = "NO";
    defparam add_1207_11.INJECT1_1 = "NO";
    CCU2D add_1207_9 (.A0(n1322[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1322[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18327), 
          .COUT(n18328), .S0(n2293[7]), .S1(n2293[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1207_9.INIT0 = 16'hf555;
    defparam add_1207_9.INIT1 = 16'hf555;
    defparam add_1207_9.INJECT1_0 = "NO";
    defparam add_1207_9.INJECT1_1 = "NO";
    CCU2D add_1207_7 (.A0(n1322[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1322[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18326), 
          .COUT(n18327), .S0(n2293[5]), .S1(n2293[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1207_7.INIT0 = 16'hf555;
    defparam add_1207_7.INIT1 = 16'hf555;
    defparam add_1207_7.INJECT1_0 = "NO";
    defparam add_1207_7.INJECT1_1 = "NO";
    CCU2D add_15135_14 (.A0(speed_set_m1[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18443), .COUT(n18444));
    defparam add_15135_14.INIT0 = 16'h5555;
    defparam add_15135_14.INIT1 = 16'h5aaa;
    defparam add_15135_14.INJECT1_0 = "NO";
    defparam add_15135_14.INJECT1_1 = "NO";
    CCU2D add_219_9 (.A0(Out2[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18261), 
          .COUT(n18262), .S0(n1343[7]), .S1(n1343[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_9.INIT0 = 16'h5aaa;
    defparam add_219_9.INIT1 = 16'h5aaa;
    defparam add_219_9.INJECT1_0 = "NO";
    defparam add_219_9.INJECT1_1 = "NO";
    CCU2D add_219_7 (.A0(Out2[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18260), 
          .COUT(n18261), .S0(n1343[5]), .S1(n1343[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_7.INIT0 = 16'h5aaa;
    defparam add_219_7.INIT1 = 16'h5aaa;
    defparam add_219_7.INJECT1_0 = "NO";
    defparam add_219_7.INJECT1_1 = "NO";
    LUT4 mux_1277_i15_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[14]), 
         .D(speed_set_m4[14]), .Z(n2613[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i15_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i4_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[3]), 
         .D(intgOut2[3]), .Z(n648[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1221_i10_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[9]), 
         .D(speed_set_m4[9]), .Z(n5407)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_138_i25_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[24]), 
         .D(intgOut2[24]), .Z(n648[24])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i12_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[11]), 
         .D(speed_set_m4[11]), .Z(n2613[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i12_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i13_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[12]), 
         .D(speed_set_m4[12]), .Z(n2613[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i13_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i12_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[11]), 
         .D(intgOut2[11]), .Z(n648[11])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i12_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i13_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[12]), 
         .D(intgOut2[12]), .Z(n648[12])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i13_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_219_5 (.A0(Out2[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18259), 
          .COUT(n18260), .S0(n1343[3]), .S1(n1343[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_5.INIT0 = 16'h5aaa;
    defparam add_219_5.INIT1 = 16'h5aaa;
    defparam add_219_5.INJECT1_0 = "NO";
    defparam add_219_5.INJECT1_1 = "NO";
    CCU2D add_219_3 (.A0(Out2[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18258), 
          .COUT(n18259), .S0(n1343[1]), .S1(n1343[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_3.INIT0 = 16'h5aaa;
    defparam add_219_3.INIT1 = 16'h5aaa;
    defparam add_219_3.INJECT1_0 = "NO";
    defparam add_219_3.INJECT1_1 = "NO";
    CCU2D add_219_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out2[13]), .B1(n18757), .C1(n18758), .D1(Out2[28]), .COUT(n18258), 
          .S1(n1343[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(336[17:21])
    defparam add_219_1.INIT0 = 16'hF000;
    defparam add_219_1.INIT1 = 16'h56aa;
    defparam add_219_1.INJECT1_0 = "NO";
    defparam add_219_1.INJECT1_1 = "NO";
    LUT4 mux_1277_i16_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[15]), 
         .D(speed_set_m4[15]), .Z(n2613[15])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i16_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_1207_5 (.A0(n1322[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1322[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18325), 
          .COUT(n18326), .S0(n2293[3]), .S1(n2293[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1207_5.INIT0 = 16'hf555;
    defparam add_1207_5.INIT1 = 16'hf555;
    defparam add_1207_5.INJECT1_0 = "NO";
    defparam add_1207_5.INJECT1_1 = "NO";
    CCU2D add_1207_3 (.A0(n1322[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1322[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18324), 
          .COUT(n18325), .S0(n2293[1]), .S1(n2293[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1207_3.INIT0 = 16'hf555;
    defparam add_1207_3.INIT1 = 16'hf555;
    defparam add_1207_3.INJECT1_0 = "NO";
    defparam add_1207_3.INJECT1_1 = "NO";
    CCU2D add_1207_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1322[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18324), 
          .S1(n2293[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(355[20:29])
    defparam add_1207_1.INIT0 = 16'hF000;
    defparam add_1207_1.INIT1 = 16'h0aaa;
    defparam add_1207_1.INJECT1_0 = "NO";
    defparam add_1207_1.INJECT1_1 = "NO";
    CCU2D add_15135_12 (.A0(speed_set_m1[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18442), .COUT(n18443));
    defparam add_15135_12.INIT0 = 16'h5aaa;
    defparam add_15135_12.INIT1 = 16'h5aaa;
    defparam add_15135_12.INJECT1_0 = "NO";
    defparam add_15135_12.INJECT1_1 = "NO";
    CCU2D add_215_17 (.A0(Out1[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18257), 
          .S0(n1322[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_17.INIT0 = 16'h5aaa;
    defparam add_215_17.INIT1 = 16'h0000;
    defparam add_215_17.INJECT1_0 = "NO";
    defparam add_215_17.INJECT1_1 = "NO";
    CCU2D add_1206_5 (.A0(n1301[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1301[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18227), 
          .COUT(n18228), .S0(n2281[3]), .S1(n2281[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(347[20:29])
    defparam add_1206_5.INIT0 = 16'hf555;
    defparam add_1206_5.INIT1 = 16'hf555;
    defparam add_1206_5.INJECT1_0 = "NO";
    defparam add_1206_5.INJECT1_1 = "NO";
    CCU2D add_215_15 (.A0(Out1[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18256), 
          .COUT(n18257), .S0(n1322[13]), .S1(n1322[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_15.INIT0 = 16'h5aaa;
    defparam add_215_15.INIT1 = 16'h5aaa;
    defparam add_215_15.INJECT1_0 = "NO";
    defparam add_215_15.INJECT1_1 = "NO";
    CCU2D add_215_13 (.A0(Out1[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18255), 
          .COUT(n18256), .S0(n1322[11]), .S1(n1322[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_13.INIT0 = 16'h5aaa;
    defparam add_215_13.INIT1 = 16'h5aaa;
    defparam add_215_13.INJECT1_0 = "NO";
    defparam add_215_13.INJECT1_1 = "NO";
    CCU2D add_15135_10 (.A0(speed_set_m1[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18441), .COUT(n18442));
    defparam add_15135_10.INIT0 = 16'h5555;
    defparam add_15135_10.INIT1 = 16'h5555;
    defparam add_15135_10.INJECT1_0 = "NO";
    defparam add_15135_10.INJECT1_1 = "NO";
    LUT4 mux_138_i24_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[23]), 
         .D(intgOut2[23]), .Z(n648[23])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i24_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i10_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[9]), 
         .D(intgOut2[9]), .Z(n648[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i10_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15135_8 (.A0(speed_set_m1[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18440), .COUT(n18441));
    defparam add_15135_8.INIT0 = 16'h5aaa;
    defparam add_15135_8.INIT1 = 16'h5555;
    defparam add_15135_8.INJECT1_0 = "NO";
    defparam add_15135_8.INJECT1_1 = "NO";
    CCU2D add_15126_17 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18497), .S1(n3752));
    defparam add_15126_17.INIT0 = 16'h5555;
    defparam add_15126_17.INIT1 = 16'h0000;
    defparam add_15126_17.INJECT1_0 = "NO";
    defparam add_15126_17.INJECT1_1 = "NO";
    CCU2D add_215_11 (.A0(Out1[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18254), 
          .COUT(n18255), .S0(n1322[9]), .S1(n1322[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_11.INIT0 = 16'h5aaa;
    defparam add_215_11.INIT1 = 16'h5aaa;
    defparam add_215_11.INJECT1_0 = "NO";
    defparam add_215_11.INJECT1_1 = "NO";
    CCU2D add_15126_15 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18496), .COUT(n18497));
    defparam add_15126_15.INIT0 = 16'hf555;
    defparam add_15126_15.INIT1 = 16'hf555;
    defparam add_15126_15.INJECT1_0 = "NO";
    defparam add_15126_15.INJECT1_1 = "NO";
    CCU2D add_15135_6 (.A0(speed_set_m1[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18439), .COUT(n18440));
    defparam add_15135_6.INIT0 = 16'h5aaa;
    defparam add_15135_6.INIT1 = 16'h5aaa;
    defparam add_15135_6.INJECT1_0 = "NO";
    defparam add_15135_6.INJECT1_1 = "NO";
    CCU2D add_215_9 (.A0(Out1[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18253), 
          .COUT(n18254), .S0(n1322[7]), .S1(n1322[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_9.INIT0 = 16'h5aaa;
    defparam add_215_9.INIT1 = 16'h5aaa;
    defparam add_215_9.INJECT1_0 = "NO";
    defparam add_215_9.INJECT1_1 = "NO";
    CCU2D add_215_7 (.A0(Out1[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18252), 
          .COUT(n18253), .S0(n1322[5]), .S1(n1322[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_7.INIT0 = 16'h5aaa;
    defparam add_215_7.INIT1 = 16'h5aaa;
    defparam add_215_7.INJECT1_0 = "NO";
    defparam add_215_7.INJECT1_1 = "NO";
    CCU2D add_215_5 (.A0(Out1[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18251), 
          .COUT(n18252), .S0(n1322[3]), .S1(n1322[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_5.INIT0 = 16'h5aaa;
    defparam add_215_5.INIT1 = 16'h5aaa;
    defparam add_215_5.INJECT1_0 = "NO";
    defparam add_215_5.INJECT1_1 = "NO";
    LUT4 mux_138_i14_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[13]), 
         .D(intgOut2[13]), .Z(n648[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i14_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_215_3 (.A0(Out1[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18250), 
          .COUT(n18251), .S0(n1322[1]), .S1(n1322[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_3.INIT0 = 16'h5aaa;
    defparam add_215_3.INIT1 = 16'h5aaa;
    defparam add_215_3.INJECT1_0 = "NO";
    defparam add_215_3.INJECT1_1 = "NO";
    LUT4 mux_138_i15_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[14]), 
         .D(intgOut2[14]), .Z(n648[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i15_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15135_4 (.A0(speed_set_m1[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18438), .COUT(n18439));
    defparam add_15135_4.INIT0 = 16'h5555;
    defparam add_15135_4.INIT1 = 16'h5aaa;
    defparam add_15135_4.INJECT1_0 = "NO";
    defparam add_15135_4.INJECT1_1 = "NO";
    CCU2D add_15135_2 (.A0(speed_set_m1[1]), .B0(speed_set_m1[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18438));
    defparam add_15135_2.INIT0 = 16'h1000;
    defparam add_15135_2.INIT1 = 16'h5555;
    defparam add_15135_2.INJECT1_0 = "NO";
    defparam add_15135_2.INJECT1_1 = "NO";
    CCU2D add_15126_13 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18495), .COUT(n18496));
    defparam add_15126_13.INIT0 = 16'hf555;
    defparam add_15126_13.INIT1 = 16'hf555;
    defparam add_15126_13.INJECT1_0 = "NO";
    defparam add_15126_13.INJECT1_1 = "NO";
    CCU2D add_215_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out1[13]), .B1(n18721), .C1(n18722), .D1(Out1[28]), .COUT(n18250), 
          .S1(n1322[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(335[17:21])
    defparam add_215_1.INIT0 = 16'hF000;
    defparam add_215_1.INIT1 = 16'h56aa;
    defparam add_215_1.INJECT1_0 = "NO";
    defparam add_215_1.INJECT1_1 = "NO";
    LUT4 mux_1277_i17_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[16]), 
         .D(speed_set_m4[16]), .Z(n2613[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i17_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_211_17 (.A0(Out0[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18249), 
          .S0(n1301[15]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_17.INIT0 = 16'h5aaa;
    defparam add_211_17.INIT1 = 16'h0000;
    defparam add_211_17.INJECT1_0 = "NO";
    defparam add_211_17.INJECT1_1 = "NO";
    FD1P3IX intgOut1_i0 (.D(addOut[0]), .SP(clk_N_875_enable_359), .CD(n15130), 
            .CK(clk_N_875), .Q(intgOut1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i0.GSR = "ENABLED";
    CCU2D add_15128_17 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18437), .S1(n3704));
    defparam add_15128_17.INIT0 = 16'h5555;
    defparam add_15128_17.INIT1 = 16'h0000;
    defparam add_15128_17.INJECT1_0 = "NO";
    defparam add_15128_17.INJECT1_1 = "NO";
    CCU2D add_15128_15 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18436), .COUT(n18437));
    defparam add_15128_15.INIT0 = 16'hf555;
    defparam add_15128_15.INIT1 = 16'hf555;
    defparam add_15128_15.INJECT1_0 = "NO";
    defparam add_15128_15.INJECT1_1 = "NO";
    LUT4 mux_1277_i18_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[17]), 
         .D(speed_set_m4[17]), .Z(n2613[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i18_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15126_11 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18494), .COUT(n18495));
    defparam add_15126_11.INIT0 = 16'hf555;
    defparam add_15126_11.INIT1 = 16'hf555;
    defparam add_15126_11.INJECT1_0 = "NO";
    defparam add_15126_11.INJECT1_1 = "NO";
    LUT4 mux_1277_i19_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[18]), 
         .D(speed_set_m4[18]), .Z(n2613[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i19_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i20_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[19]), 
         .D(intgOut2[19]), .Z(n648[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i20_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1221_i7_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[6]), 
         .D(speed_set_m4[6]), .Z(n5401)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i7_3_lut_4_lut.init = 16'hf780;
    FD1P3IX intgOut0_i0 (.D(addOut[0]), .SP(clk_N_875_enable_387), .CD(n14299), 
            .CK(clk_N_875), .Q(intgOut0[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i0.GSR = "ENABLED";
    LUT4 mux_1277_i20_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[19]), 
         .D(speed_set_m4[19]), .Z(n2613[19])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i20_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i21_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[20]), 
         .D(speed_set_m4[20]), .Z(n2613[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i17_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[16]), 
         .D(intgOut2[16]), .Z(n648[16])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i17_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i18_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[17]), 
         .D(intgOut2[17]), .Z(n648[17])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i18_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i1_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[0]), 
         .D(speed_set_m4[0]), .Z(n2613[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1221_i5_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[4]), 
         .D(speed_set_m4[4]), .Z(n5397)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_138_i19_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[18]), 
         .D(intgOut2[18]), .Z(n648[18])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i19_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i23_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[22]), 
         .D(intgOut2[22]), .Z(n648[22])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i23_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i4_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[3]), 
         .D(speed_set_m4[3]), .Z(n2613[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i8_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[7]), 
         .D(speed_set_m4[7]), .Z(n2613[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i3_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[2]), 
         .D(intgOut2[2]), .Z(n648[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i9_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[8]), 
         .D(speed_set_m4[8]), .Z(n2613[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i9_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i5_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[4]), 
         .D(intgOut2[4]), .Z(n648[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i5_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i6_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[5]), 
         .D(speed_set_m4[5]), .Z(n2613[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 i14064_3_lut_4_lut (.A(n21465), .B(n21466), .C(n4_adj_2364), 
         .D(n3776), .Z(n16674)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i14064_3_lut_4_lut.init = 16'hfeee;
    LUT4 mux_1277_i10_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[9]), 
         .D(speed_set_m4[9]), .Z(n2613[9])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i10_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15128_13 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18435), .COUT(n18436));
    defparam add_15128_13.INIT0 = 16'hf555;
    defparam add_15128_13.INIT1 = 16'hf555;
    defparam add_15128_13.INJECT1_0 = "NO";
    defparam add_15128_13.INJECT1_1 = "NO";
    LUT4 mux_1222_i8_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[7]), 
         .D(speed_set_m3[7]), .Z(n5361)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1221_i4_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[3]), 
         .D(speed_set_m4[3]), .Z(n5395)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1277_i11_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[10]), 
         .D(speed_set_m4[10]), .Z(n2613[10])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i11_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i6_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[5]), 
         .D(intgOut2[5]), .Z(n648[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i7_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[6]), 
         .D(intgOut2[6]), .Z(n648[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i3_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[2]), 
         .D(speed_set_m4[2]), .Z(n2613[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13415_2_lut (.A(addOut[16]), .B(n22216), .Z(backOut3_28__N_1874[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13415_2_lut.init = 16'h2222;
    LUT4 mux_1277_i14_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[13]), 
         .D(speed_set_m4[13]), .Z(n2613[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i14_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i28_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[27]), 
         .D(intgOut2[27]), .Z(n648[27])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i28_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_15128_11 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18434), .COUT(n18435));
    defparam add_15128_11.INIT0 = 16'hf555;
    defparam add_15128_11.INIT1 = 16'hf555;
    defparam add_15128_11.INJECT1_0 = "NO";
    defparam add_15128_11.INJECT1_1 = "NO";
    CCU2D add_15128_9 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18433), .COUT(n18434));
    defparam add_15128_9.INIT0 = 16'hf555;
    defparam add_15128_9.INIT1 = 16'h0aaa;
    defparam add_15128_9.INJECT1_0 = "NO";
    defparam add_15128_9.INJECT1_1 = "NO";
    CCU2D add_15126_9 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18493), .COUT(n18494));
    defparam add_15126_9.INIT0 = 16'hf555;
    defparam add_15126_9.INIT1 = 16'h0aaa;
    defparam add_15126_9.INJECT1_0 = "NO";
    defparam add_15126_9.INJECT1_1 = "NO";
    LUT4 mux_138_i8_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[7]), 
         .D(intgOut2[7]), .Z(n648[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i5_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[4]), 
         .D(speed_set_m4[4]), .Z(n2613[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i5_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i29_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[28]), 
         .D(intgOut2[28]), .Z(n648[28])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i29_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1221_i15_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[14]), 
         .D(speed_set_m4[14]), .Z(n5417)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_138_i9_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[8]), 
         .D(intgOut2[8]), .Z(n648[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i9_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_138_i21_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[20]), 
         .D(intgOut2[20]), .Z(n648[20])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i21_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1277_i7_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[6]), 
         .D(speed_set_m4[6]), .Z(n2613[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 i13414_2_lut (.A(addOut[15]), .B(n22216), .Z(backOut3_28__N_1874[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13414_2_lut.init = 16'h2222;
    LUT4 mux_1277_i2_3_lut_4_lut (.A(n15773), .B(n49), .C(speed_set_m3[1]), 
         .D(speed_set_m4[1]), .Z(n2613[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_1277_i2_3_lut_4_lut.init = 16'hfe10;
    LUT4 ss_3__bdd_4_lut (.A(ss[3]), .B(n6), .C(n21444), .D(n22216), 
         .Z(n15757)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam ss_3__bdd_4_lut.init = 16'hf0d0;
    LUT4 i1_2_lut_adj_116 (.A(ss[0]), .B(ss[3]), .Z(n11644)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_adj_116.init = 16'h8888;
    LUT4 n9_bdd_4_lut (.A(n21443), .B(n21467), .C(ss[0]), .D(ss[1]), 
         .Z(n15773)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))) */ ;
    defparam n9_bdd_4_lut.init = 16'ha88a;
    LUT4 mux_1221_i20_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[19]), 
         .D(speed_set_m4[19]), .Z(n5427)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_138_i1_3_lut_4_lut (.A(n21465), .B(n21467), .C(intgOut1[0]), 
         .D(intgOut2[0]), .Z(n648[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(169[9:16])
    defparam mux_138_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_adj_117 (.A(n1364[15]), .B(n2317[9]), .C(n30_adj_2374), 
         .Z(n19131)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[4] 376[11])
    defparam i1_3_lut_adj_117.init = 16'h8a8a;
    CCU2D add_211_15 (.A0(Out0[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18248), 
          .COUT(n18249), .S0(n1301[13]), .S1(n1301[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_15.INIT0 = 16'h5aaa;
    defparam add_211_15.INIT1 = 16'h5aaa;
    defparam add_211_15.INJECT1_0 = "NO";
    defparam add_211_15.INJECT1_1 = "NO";
    LUT4 i5_4_lut_adj_118 (.A(n9_adj_2375), .B(n7), .C(n1364[10]), .D(n1364[13]), 
         .Z(n30_adj_2374)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_118.init = 16'h8000;
    CCU2D add_15126_7 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18492), .COUT(n18493));
    defparam add_15126_7.INIT0 = 16'h0aaa;
    defparam add_15126_7.INIT1 = 16'hf555;
    defparam add_15126_7.INJECT1_0 = "NO";
    defparam add_15126_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_119 (.A(n1343[15]), .B(n2305[7]), .C(n9_adj_2373), 
         .Z(n1502[7])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_119.init = 16'h8a8a;
    LUT4 i3_2_lut_adj_120 (.A(n1364[14]), .B(n1364[12]), .Z(n9_adj_2375)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_120.init = 16'h8888;
    CCU2D add_15126_5 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18491), .COUT(n18492));
    defparam add_15126_5.INIT0 = 16'h0aaa;
    defparam add_15126_5.INIT1 = 16'h0aaa;
    defparam add_15126_5.INJECT1_0 = "NO";
    defparam add_15126_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_121 (.A(n1364[11]), .B(n1364[9]), .C(n10_adj_2376), 
         .D(n1364[7]), .Z(n7)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_121.init = 16'haaa8;
    LUT4 i4_4_lut_adj_122 (.A(n1364[6]), .B(n8_adj_2377), .C(n1364[4]), 
         .D(n4_adj_2378), .Z(n10_adj_2376)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_122.init = 16'hfeee;
    LUT4 i2_2_lut_adj_123 (.A(n1364[5]), .B(n1364[8]), .Z(n8_adj_2377)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_123.init = 16'heeee;
    LUT4 i1_4_lut_adj_124 (.A(n1364[3]), .B(n1364[2]), .C(n1364[1]), .D(n1364[0]), 
         .Z(n4_adj_2378)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_124.init = 16'haaa8;
    LUT4 i1_3_lut_adj_125 (.A(n1364[15]), .B(n2317[8]), .C(n30_adj_2374), 
         .Z(n19125)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[4] 376[11])
    defparam i1_3_lut_adj_125.init = 16'h8a8a;
    LUT4 i13413_2_lut (.A(addOut[14]), .B(n22216), .Z(backOut3_28__N_1874[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13413_2_lut.init = 16'h2222;
    LUT4 i52_2_lut_rep_307 (.A(n15773), .B(n49), .Z(n21408)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(138[23] 139[51])
    defparam i52_2_lut_rep_307.init = 16'h4444;
    LUT4 i13412_2_lut (.A(addOut[13]), .B(n22216), .Z(backOut3_28__N_1874[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13412_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_adj_126 (.A(n15773), .B(n49), .C(n11585), .D(n21409), 
         .Z(n2565)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(138[23] 139[51])
    defparam i1_3_lut_4_lut_adj_126.init = 16'hf040;
    LUT4 i1_3_lut_adj_127 (.A(n1364[15]), .B(n2317[7]), .C(n30_adj_2374), 
         .Z(n19119)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(370[4] 376[11])
    defparam i1_3_lut_adj_127.init = 16'h8a8a;
    LUT4 i1_3_lut_adj_128 (.A(n1364[15]), .B(n2317[6]), .C(n30_adj_2374), 
         .Z(n1546[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_128.init = 16'h8a8a;
    LUT4 i1_2_lut_rep_308 (.A(n16496), .B(n42), .Z(n21409)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam i1_2_lut_rep_308.init = 16'h4444;
    LUT4 mux_1222_i5_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[4]), 
         .D(speed_set_m3[4]), .Z(n5355)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1222_i14_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[13]), 
         .D(speed_set_m3[13]), .Z(n5373)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1222_i21_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[20]), 
         .D(speed_set_m3[20]), .Z(n5387)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_adj_129 (.A(n1364[15]), .B(n2317[5]), .C(n30_adj_2374), 
         .Z(n1546[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_129.init = 16'h8a8a;
    LUT4 mux_1222_i19_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[18]), 
         .D(speed_set_m3[18]), .Z(n5383)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1221_i21_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[20]), 
         .D(speed_set_m4[20]), .Z(n5429)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1222_i18_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[17]), 
         .D(speed_set_m3[17]), .Z(n5381)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13411_2_lut (.A(addOut[12]), .B(n22216), .Z(backOut3_28__N_1874[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13411_2_lut.init = 16'h2222;
    LUT4 mux_1222_i9_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[8]), 
         .D(speed_set_m3[8]), .Z(n5363)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1222_i4_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[3]), 
         .D(speed_set_m3[3]), .Z(n5353)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_1222_i13_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[12]), 
         .D(speed_set_m3[12]), .Z(n5371)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13601_2_lut (.A(addOut[11]), .B(n22216), .Z(Out2_28__N_1145[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13601_2_lut.init = 16'h2222;
    LUT4 i13407_2_lut (.A(addOut[10]), .B(n22216), .Z(backOut3_28__N_1874[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13407_2_lut.init = 16'h2222;
    PFUMX mux_1226_i21 (.BLUT(n5429), .ALUT(n5387), .C0(n2565), .Z(n5473));
    PFUMX mux_1226_i20 (.BLUT(n5427), .ALUT(n5385), .C0(n2565), .Z(n5471));
    PFUMX mux_1226_i19 (.BLUT(n5425), .ALUT(n5383), .C0(n2565), .Z(n5469));
    PFUMX mux_1226_i18 (.BLUT(n5423), .ALUT(n5381), .C0(n2565), .Z(n5467));
    LUT4 mux_1222_i20_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[19]), 
         .D(speed_set_m3[19]), .Z(n5385)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 i13406_2_lut (.A(addOut[9]), .B(n22216), .Z(backOut3_28__N_1874[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13406_2_lut.init = 16'h2222;
    LUT4 i13405_2_lut (.A(addOut[8]), .B(n22216), .Z(backOut3_28__N_1874[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13405_2_lut.init = 16'h2222;
    PFUMX mux_1226_i17 (.BLUT(n5421), .ALUT(n5379), .C0(n2565), .Z(n5465));
    LUT4 i13400_2_lut (.A(addOut[7]), .B(n22216), .Z(backOut3_28__N_1874[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13400_2_lut.init = 16'h2222;
    LUT4 i13393_2_lut (.A(addOut[6]), .B(n22216), .Z(backOut3_28__N_1874[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13393_2_lut.init = 16'h2222;
    LUT4 i11833_4_lut (.A(clk_N_875_enable_391), .B(n21463), .C(n30_adj_2374), 
         .D(n1364[15]), .Z(n14437)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11833_4_lut.init = 16'h8aaa;
    PFUMX mux_1226_i16 (.BLUT(n5419), .ALUT(n5377), .C0(n2565), .Z(n5463));
    PFUMX mux_1226_i15 (.BLUT(n5417), .ALUT(n5375), .C0(n2565), .Z(n5461));
    LUT4 i1_3_lut_adj_130 (.A(n1364[15]), .B(n2317[3]), .C(n30_adj_2374), 
         .Z(n1546[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_130.init = 16'h8a8a;
    PFUMX mux_1226_i14 (.BLUT(n5415), .ALUT(n5373), .C0(n2565), .Z(n5459));
    PFUMX mux_1226_i13 (.BLUT(n5413), .ALUT(n5371), .C0(n2565), .Z(n5457));
    LUT4 i13384_2_lut (.A(addOut[5]), .B(n22216), .Z(backOut3_28__N_1874[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13384_2_lut.init = 16'h2222;
    CCU2D add_15128_7 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18432), .COUT(n18433));
    defparam add_15128_7.INIT0 = 16'h0aaa;
    defparam add_15128_7.INIT1 = 16'hf555;
    defparam add_15128_7.INJECT1_0 = "NO";
    defparam add_15128_7.INJECT1_1 = "NO";
    CCU2D add_211_13 (.A0(Out0[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18247), 
          .COUT(n18248), .S0(n1301[11]), .S1(n1301[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_13.INIT0 = 16'h5aaa;
    defparam add_211_13.INIT1 = 16'h5aaa;
    defparam add_211_13.INJECT1_0 = "NO";
    defparam add_211_13.INJECT1_1 = "NO";
    PFUMX mux_1226_i12 (.BLUT(n5411), .ALUT(n5369), .C0(n2565), .Z(n5455));
    PFUMX mux_1226_i11 (.BLUT(n5409), .ALUT(n5367), .C0(n2565), .Z(n5453));
    CCU2D add_211_11 (.A0(Out0[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18246), 
          .COUT(n18247), .S0(n1301[9]), .S1(n1301[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_11.INIT0 = 16'h5aaa;
    defparam add_211_11.INIT1 = 16'h5aaa;
    defparam add_211_11.INJECT1_0 = "NO";
    defparam add_211_11.INJECT1_1 = "NO";
    PFUMX mux_1226_i10 (.BLUT(n5407), .ALUT(n5365), .C0(n2565), .Z(n5451));
    PFUMX mux_1226_i9 (.BLUT(n5405), .ALUT(n5363), .C0(n2565), .Z(n5449));
    PFUMX mux_1226_i8 (.BLUT(n5403), .ALUT(n5361), .C0(n2565), .Z(n5447));
    PFUMX mux_1226_i7 (.BLUT(n5401), .ALUT(n5359), .C0(n2565), .Z(n5445));
    CCU2D add_15128_5 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18431), .COUT(n18432));
    defparam add_15128_5.INIT0 = 16'h0aaa;
    defparam add_15128_5.INIT1 = 16'h0aaa;
    defparam add_15128_5.INJECT1_0 = "NO";
    defparam add_15128_5.INJECT1_1 = "NO";
    CCU2D add_15128_3 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18430), .COUT(n18431));
    defparam add_15128_3.INIT0 = 16'hf555;
    defparam add_15128_3.INIT1 = 16'hf555;
    defparam add_15128_3.INJECT1_0 = "NO";
    defparam add_15128_3.INJECT1_1 = "NO";
    CCU2D add_15128_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[4]), .B1(speed_set_m3[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18430));
    defparam add_15128_1.INIT0 = 16'hF000;
    defparam add_15128_1.INIT1 = 16'ha666;
    defparam add_15128_1.INJECT1_0 = "NO";
    defparam add_15128_1.INJECT1_1 = "NO";
    PFUMX mux_1226_i6 (.BLUT(n5399), .ALUT(n5357), .C0(n2565), .Z(n5443));
    LUT4 i13383_2_lut (.A(addOut[4]), .B(n22216), .Z(backOut3_28__N_1874[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13383_2_lut.init = 16'h2222;
    PFUMX mux_1226_i5 (.BLUT(n5397), .ALUT(n5355), .C0(n2565), .Z(n5441));
    LUT4 i13382_2_lut (.A(addOut[3]), .B(n22216), .Z(backOut3_28__N_1874[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13382_2_lut.init = 16'h2222;
    CCU2D add_15126_3 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18490), .COUT(n18491));
    defparam add_15126_3.INIT0 = 16'hf555;
    defparam add_15126_3.INIT1 = 16'hf555;
    defparam add_15126_3.INJECT1_0 = "NO";
    defparam add_15126_3.INJECT1_1 = "NO";
    LUT4 i13381_2_lut (.A(addOut[2]), .B(n22216), .Z(backOut3_28__N_1874[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13381_2_lut.init = 16'h2222;
    CCU2D add_15126_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[4]), .B1(speed_set_m4[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18490));
    defparam add_15126_1.INIT0 = 16'hF000;
    defparam add_15126_1.INIT1 = 16'ha666;
    defparam add_15126_1.INJECT1_0 = "NO";
    defparam add_15126_1.INJECT1_1 = "NO";
    CCU2D add_211_9 (.A0(Out0[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18245), 
          .COUT(n18246), .S0(n1301[7]), .S1(n1301[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_9.INIT0 = 16'h5aaa;
    defparam add_211_9.INIT1 = 16'h5aaa;
    defparam add_211_9.INJECT1_0 = "NO";
    defparam add_211_9.INJECT1_1 = "NO";
    LUT4 i13378_2_lut (.A(addOut[1]), .B(n22216), .Z(backOut3_28__N_1874[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i13378_2_lut.init = 16'h2222;
    PFUMX mux_1226_i4 (.BLUT(n5395), .ALUT(n5353), .C0(n2565), .Z(n5439));
    PFUMX mux_1226_i3 (.BLUT(n5393), .ALUT(n5351), .C0(n2565), .Z(n5437));
    CCU2D add_15129_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18303), 
          .S0(n3776));
    defparam add_15129_cout.INIT0 = 16'h0000;
    defparam add_15129_cout.INIT1 = 16'h0000;
    defparam add_15129_cout.INJECT1_0 = "NO";
    defparam add_15129_cout.INJECT1_1 = "NO";
    PFUMX mux_1226_i2 (.BLUT(n5391), .ALUT(n5349), .C0(n2565), .Z(n5435));
    CCU2D add_15129_20 (.A0(speed_set_m4[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18302), .COUT(n18303));
    defparam add_15129_20.INIT0 = 16'h5aaa;
    defparam add_15129_20.INIT1 = 16'h0aaa;
    defparam add_15129_20.INJECT1_0 = "NO";
    defparam add_15129_20.INJECT1_1 = "NO";
    LUT4 i3_2_lut_adj_131 (.A(n1322[14]), .B(n1322[12]), .Z(n9_adj_2379)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_131.init = 16'h8888;
    PFUMX mux_1226_i1 (.BLUT(n5347), .ALUT(n5345), .C0(n2565), .Z(n5433));
    PFUMX i3055 (.BLUT(n2613[0]), .ALUT(n5556), .C0(n21403), .Z(n5557));
    PFUMX i3367 (.BLUT(n2613[1]), .ALUT(n5868), .C0(n21403), .Z(n5869));
    PFUMX i3369 (.BLUT(n2613[2]), .ALUT(n5870), .C0(n21403), .Z(n5871));
    PFUMX i3371 (.BLUT(n2613[3]), .ALUT(n5872), .C0(n21403), .Z(n5873));
    PFUMX i3373 (.BLUT(n2613[4]), .ALUT(n5874), .C0(n21403), .Z(n5875));
    CCU2D add_15129_18 (.A0(speed_set_m4[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18301), .COUT(n18302));
    defparam add_15129_18.INIT0 = 16'h5aaa;
    defparam add_15129_18.INIT1 = 16'h5aaa;
    defparam add_15129_18.INJECT1_0 = "NO";
    defparam add_15129_18.INJECT1_1 = "NO";
    CCU2D add_15129_16 (.A0(speed_set_m4[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18300), .COUT(n18301));
    defparam add_15129_16.INIT0 = 16'h5aaa;
    defparam add_15129_16.INIT1 = 16'h5aaa;
    defparam add_15129_16.INJECT1_0 = "NO";
    defparam add_15129_16.INJECT1_1 = "NO";
    CCU2D add_211_7 (.A0(Out0[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18244), 
          .COUT(n18245), .S0(n1301[5]), .S1(n1301[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_7.INIT0 = 16'h5aaa;
    defparam add_211_7.INIT1 = 16'h5aaa;
    defparam add_211_7.INJECT1_0 = "NO";
    defparam add_211_7.INJECT1_1 = "NO";
    PFUMX i3375 (.BLUT(n2613[5]), .ALUT(n5876), .C0(n21403), .Z(n5877));
    PFUMX i3377 (.BLUT(n2613[6]), .ALUT(n5878), .C0(n21403), .Z(n5879));
    PFUMX i3379 (.BLUT(n2613[7]), .ALUT(n5880), .C0(n21403), .Z(n5881));
    PFUMX i3381 (.BLUT(n2613[8]), .ALUT(n5882), .C0(n21403), .Z(n5883));
    PFUMX i3383 (.BLUT(n2613[9]), .ALUT(n5884), .C0(n21403), .Z(n5885));
    LUT4 i1_3_lut_adj_132 (.A(n1343[15]), .B(n2305[9]), .C(n9_adj_2373), 
         .Z(n1502[9])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_132.init = 16'h8a8a;
    PFUMX i3385 (.BLUT(n2613[10]), .ALUT(n5886), .C0(n21403), .Z(n5887));
    PFUMX i3387 (.BLUT(n2613[11]), .ALUT(n5888), .C0(n21403), .Z(n5889));
    PFUMX i3389 (.BLUT(n2613[12]), .ALUT(n5890), .C0(n21403), .Z(n5891));
    PFUMX i3391 (.BLUT(n2613[13]), .ALUT(n5892), .C0(n21403), .Z(n5893));
    PFUMX i3393 (.BLUT(n2613[14]), .ALUT(n5894), .C0(n21403), .Z(n5895));
    CCU2D add_15129_14 (.A0(speed_set_m4[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18299), .COUT(n18300));
    defparam add_15129_14.INIT0 = 16'h5555;
    defparam add_15129_14.INIT1 = 16'h5aaa;
    defparam add_15129_14.INJECT1_0 = "NO";
    defparam add_15129_14.INJECT1_1 = "NO";
    CCU2D add_15129_12 (.A0(speed_set_m4[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18298), .COUT(n18299));
    defparam add_15129_12.INIT0 = 16'h5aaa;
    defparam add_15129_12.INIT1 = 16'h5aaa;
    defparam add_15129_12.INJECT1_0 = "NO";
    defparam add_15129_12.INJECT1_1 = "NO";
    CCU2D add_15129_10 (.A0(speed_set_m4[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18297), .COUT(n18298));
    defparam add_15129_10.INIT0 = 16'h5555;
    defparam add_15129_10.INIT1 = 16'h5555;
    defparam add_15129_10.INJECT1_0 = "NO";
    defparam add_15129_10.INJECT1_1 = "NO";
    CCU2D add_211_5 (.A0(Out0[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18243), 
          .COUT(n18244), .S0(n1301[3]), .S1(n1301[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_5.INIT0 = 16'h5aaa;
    defparam add_211_5.INIT1 = 16'h5aaa;
    defparam add_211_5.INJECT1_0 = "NO";
    defparam add_211_5.INJECT1_1 = "NO";
    PFUMX i3395 (.BLUT(n2613[15]), .ALUT(n5896), .C0(n21403), .Z(n5897));
    PFUMX i3397 (.BLUT(n2613[16]), .ALUT(n5898), .C0(n21403), .Z(n5899));
    PFUMX i3399 (.BLUT(n2613[17]), .ALUT(n5900), .C0(n21403), .Z(n5901));
    LUT4 i5_4_lut_adj_133 (.A(n9_adj_2380), .B(n1343[10]), .C(n8_adj_2381), 
         .D(n1343[11]), .Z(n9_adj_2373)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_133.init = 16'h8000;
    PFUMX i3401 (.BLUT(n2613[18]), .ALUT(n5902), .C0(n21403), .Z(n5903));
    PFUMX i3403 (.BLUT(n2613[19]), .ALUT(n5904), .C0(n21403), .Z(n5905));
    PFUMX i3407 (.BLUT(n2613[20]), .ALUT(n5908), .C0(n21403), .Z(n5909));
    CCU2D add_15129_8 (.A0(speed_set_m4[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18296), .COUT(n18297));
    defparam add_15129_8.INIT0 = 16'h5aaa;
    defparam add_15129_8.INIT1 = 16'h5555;
    defparam add_15129_8.INJECT1_0 = "NO";
    defparam add_15129_8.INJECT1_1 = "NO";
    LUT4 i3_2_lut_adj_134 (.A(n1343[14]), .B(n1343[13]), .Z(n9_adj_2380)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut_adj_134.init = 16'h8888;
    L6MUX21 addIn2_28__I_29_i14 (.D0(n618[13]), .D1(addIn2_28__N_1571[13]), 
            .SD(n20127), .Z(addIn2_28__N_1441[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i15 (.D0(n618[14]), .D1(addIn2_28__N_1571[14]), 
            .SD(n20127), .Z(addIn2_28__N_1441[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i16 (.D0(n618[15]), .D1(addIn2_28__N_1571[15]), 
            .SD(n20127), .Z(addIn2_28__N_1441[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i17 (.D0(n618[16]), .D1(addIn2_28__N_1571[16]), 
            .SD(n20127), .Z(addIn2_28__N_1441[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i18 (.D0(n618[17]), .D1(addIn2_28__N_1571[17]), 
            .SD(n20127), .Z(addIn2_28__N_1441[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i19 (.D0(n618[18]), .D1(addIn2_28__N_1571[18]), 
            .SD(n20127), .Z(addIn2_28__N_1441[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i20 (.D0(n618[19]), .D1(addIn2_28__N_1571[19]), 
            .SD(n20127), .Z(addIn2_28__N_1441[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i21 (.D0(n618[20]), .D1(addIn2_28__N_1571[20]), 
            .SD(n20127), .Z(addIn2_28__N_1441[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i2_4_lut_adj_135 (.A(n1343[9]), .B(n1343[12]), .C(n10_adj_2382), 
         .D(n1343[7]), .Z(n8_adj_2381)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_135.init = 16'hccc8;
    L6MUX21 addIn2_28__I_29_i2 (.D0(n618[1]), .D1(addIn2_28__N_1571[1]), 
            .SD(n20127), .Z(addIn2_28__N_1441[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i22 (.D0(n618[21]), .D1(addIn2_28__N_1571[21]), 
            .SD(n20127), .Z(addIn2_28__N_1441[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i4_4_lut_adj_136 (.A(n1343[6]), .B(n8_adj_2383), .C(n1343[4]), 
         .D(n4_adj_2384), .Z(n10_adj_2382)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_136.init = 16'hfeee;
    L6MUX21 addIn2_28__I_29_i3 (.D0(n618[2]), .D1(addIn2_28__N_1571[2]), 
            .SD(n20127), .Z(addIn2_28__N_1441[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i23 (.D0(n618[22]), .D1(addIn2_28__N_1571[22]), 
            .SD(n20127), .Z(addIn2_28__N_1441[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i4 (.D0(n618[3]), .D1(addIn2_28__N_1571[3]), 
            .SD(n20127), .Z(addIn2_28__N_1441[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i5 (.D0(n618[4]), .D1(addIn2_28__N_1571[4]), 
            .SD(n20127), .Z(addIn2_28__N_1441[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15133_21 (.A0(speed_set_m4[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18489), .S1(n56));
    defparam add_15133_21.INIT0 = 16'h5555;
    defparam add_15133_21.INIT1 = 16'h0000;
    defparam add_15133_21.INJECT1_0 = "NO";
    defparam add_15133_21.INJECT1_1 = "NO";
    L6MUX21 addIn2_28__I_29_i24 (.D0(n618[23]), .D1(addIn2_28__N_1571[23]), 
            .SD(n20127), .Z(addIn2_28__N_1441[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i6 (.D0(n618[5]), .D1(addIn2_28__N_1571[5]), 
            .SD(n20127), .Z(addIn2_28__N_1441[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i25 (.D0(n618[24]), .D1(addIn2_28__N_1571[24]), 
            .SD(n20127), .Z(addIn2_28__N_1441[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i7 (.D0(n618[6]), .D1(addIn2_28__N_1571[6]), 
            .SD(n20127), .Z(addIn2_28__N_1441[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i26 (.D0(n618[25]), .D1(addIn2_28__N_1571[25]), 
            .SD(n20127), .Z(addIn2_28__N_1441[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i8 (.D0(n618[7]), .D1(addIn2_28__N_1571[7]), 
            .SD(n20127), .Z(addIn2_28__N_1441[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    L6MUX21 addIn2_28__I_29_i27 (.D0(n618[26]), .D1(addIn2_28__N_1571[26]), 
            .SD(n20127), .Z(addIn2_28__N_1441[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m4_i0_i9 (.D(n19131), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m4[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i8 (.D(n19125), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m4[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i7 (.D(n19119), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m4[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i7.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i9 (.D0(n618[8]), .D1(addIn2_28__N_1571[8]), 
            .SD(n20127), .Z(addIn2_28__N_1441[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m4_i0_i6 (.D(n1546[6]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m4[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i6.GSR = "DISABLED";
    CCU2D add_15133_19 (.A0(speed_set_m4[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18488), .COUT(n18489));
    defparam add_15133_19.INIT0 = 16'hf555;
    defparam add_15133_19.INIT1 = 16'hf555;
    defparam add_15133_19.INJECT1_0 = "NO";
    defparam add_15133_19.INJECT1_1 = "NO";
    FD1P3IX dutyout_m4_i0_i5 (.D(n1546[5]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m4[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i5.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i10 (.D0(n618[9]), .D1(addIn2_28__N_1571[9]), 
            .SD(n20127), .Z(addIn2_28__N_1441[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m4_i0_i4 (.D(n2317[4]), .SP(clk_N_875_enable_391), .CD(n14437), 
            .CK(clk_N_875), .Q(PWMdut_m4[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i3 (.D(n1546[3]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m4[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i3.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i28 (.D0(n618[27]), .D1(addIn2_28__N_1571[27]), 
            .SD(n20127), .Z(addIn2_28__N_1441[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m4_i0_i2 (.D(n2317[2]), .SP(clk_N_875_enable_391), .CD(n14437), 
            .CK(clk_N_875), .Q(PWMdut_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m4_i0_i1 (.D(n2317[1]), .SP(clk_N_875_enable_391), .CD(n14437), 
            .CK(clk_N_875), .Q(PWMdut_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i9 (.D(n1502[9]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i8 (.D(n1502[8]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i8.GSR = "DISABLED";
    LUT4 mux_1221_i19_3_lut_4_lut (.A(subIn1_24__N_1342), .B(n35), .C(speed_set_m1[18]), 
         .D(speed_set_m4[18]), .Z(n5425)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(134[23] 135[50])
    defparam mux_1221_i19_3_lut_4_lut.init = 16'hf780;
    FD1P3IX dutyout_m3_i0_i7 (.D(n1502[7]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i6 (.D(n1502[6]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i5 (.D(n1502[5]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i5.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i29 (.D0(n618[28]), .D1(addIn2_28__N_1571[28]), 
            .SD(n20127), .Z(addIn2_28__N_1441[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m3_i0_i4 (.D(n2305[4]), .SP(clk_N_875_enable_391), .CD(n14428), 
            .CK(clk_N_875), .Q(PWMdut_m3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i3 (.D(n1502[3]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i2 (.D(n2305[2]), .SP(clk_N_875_enable_391), .CD(n14428), 
            .CK(clk_N_875), .Q(PWMdut_m3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i1 (.D(n2305[1]), .SP(clk_N_875_enable_391), .CD(n14428), 
            .CK(clk_N_875), .Q(PWMdut_m3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i1.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i11 (.D0(n618[10]), .D1(addIn2_28__N_1571[10]), 
            .SD(n20127), .Z(addIn2_28__N_1441[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m2_i0_i9 (.D(n19113), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i8 (.D(n19107), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i7 (.D(n19101), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i7.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i6 (.D(n1458[6]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i5 (.D(n1458[5]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i4 (.D(n2293[4]), .SP(clk_N_875_enable_391), .CD(n14419), 
            .CK(clk_N_875), .Q(PWMdut_m2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i4.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i3 (.D(n1458[3]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i2 (.D(n2293[2]), .SP(clk_N_875_enable_391), .CD(n14419), 
            .CK(clk_N_875), .Q(PWMdut_m2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i2.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i12 (.D0(n618[11]), .D1(addIn2_28__N_1571[11]), 
            .SD(n20127), .Z(addIn2_28__N_1441[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m2_i0_i1 (.D(n2293[1]), .SP(clk_N_875_enable_391), .CD(n14419), 
            .CK(clk_N_875), .Q(PWMdut_m2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i1.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i9 (.D(n1414[9]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i9.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i8 (.D(n1414[8]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i8.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i7 (.D(n1414[7]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i7.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i13 (.D0(n618[12]), .D1(addIn2_28__N_1571[12]), 
            .SD(n20127), .Z(addIn2_28__N_1441[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m1_i0_i6 (.D(n1414[6]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i6.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i5 (.D(n1414[5]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i5.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i4 (.D(n2281[4]), .SP(clk_N_875_enable_391), .CD(n14410), 
            .CK(clk_N_875), .Q(PWMdut_m1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i4.GSR = "DISABLED";
    L6MUX21 addIn2_28__I_29_i1 (.D0(n618[0]), .D1(addIn2_28__N_1571[0]), 
            .SD(n20127), .Z(addIn2_28__N_1441[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m1_i0_i3 (.D(n1414[3]), .SP(clk_N_875_enable_391), .CD(n14414), 
            .CK(clk_N_875), .Q(PWMdut_m1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i3.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i2 (.D(n2281[2]), .SP(clk_N_875_enable_391), .CD(n14410), 
            .CK(clk_N_875), .Q(PWMdut_m1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i2.GSR = "DISABLED";
    FD1P3IX dutyout_m1_i0_i1 (.D(n2281[1]), .SP(clk_N_875_enable_391), .CD(n14410), 
            .CK(clk_N_875), .Q(PWMdut_m1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i1.GSR = "DISABLED";
    FD1P3IX intgOut3_i28 (.D(intgOut0_28__N_1629[28]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i28.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i13 (.BLUT(n367[12]), .ALUT(subIn2_24__N_1348[12]), 
          .C0(n20374), .Z(n4447)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i27 (.D(intgOut0_28__N_1629[27]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i27.GSR = "ENABLED";
    FD1P3IX intgOut3_i26 (.D(intgOut0_28__N_1629[26]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i26.GSR = "ENABLED";
    FD1P3IX intgOut3_i25 (.D(intgOut0_28__N_1629[25]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i25.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i10 (.BLUT(n367[9]), .ALUT(subIn2_24__N_1348[9]), 
          .C0(n20374), .Z(n4450)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i24 (.D(intgOut0_28__N_1629[24]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i24.GSR = "ENABLED";
    FD1P3IX intgOut3_i23 (.D(intgOut0_28__N_1629[23]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i23.GSR = "ENABLED";
    FD1P3IX intgOut3_i22 (.D(intgOut0_28__N_1629[22]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i22.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i9 (.BLUT(n367[8]), .ALUT(subIn2_24__N_1348[8]), 
          .C0(n20374), .Z(n4451)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i21 (.D(intgOut0_28__N_1629[21]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i21.GSR = "ENABLED";
    CCU2D add_15133_17 (.A0(speed_set_m4[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18487), .COUT(n18488));
    defparam add_15133_17.INIT0 = 16'hf555;
    defparam add_15133_17.INIT1 = 16'hf555;
    defparam add_15133_17.INJECT1_0 = "NO";
    defparam add_15133_17.INJECT1_1 = "NO";
    PFUMX subIn2_24__I_0_rep_1_i8 (.BLUT(n367[7]), .ALUT(subIn2_24__N_1348[7]), 
          .C0(n20374), .Z(n4452)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i20 (.D(intgOut0_28__N_1629[20]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i20.GSR = "ENABLED";
    FD1P3IX intgOut3_i19 (.D(intgOut0_28__N_1629[19]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i19.GSR = "ENABLED";
    FD1P3IX intgOut3_i18 (.D(intgOut0_28__N_1629[18]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i18.GSR = "ENABLED";
    FD1P3IX intgOut3_i17 (.D(intgOut0_28__N_1629[17]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i17.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i4 (.BLUT(n367[3]), .ALUT(subIn2_24__N_1348[3]), 
          .C0(n20374), .Z(n4456)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i16 (.D(intgOut0_28__N_1629[16]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i16.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i20 (.BLUT(subIn2_24__N_1535[19]), .ALUT(subIn2_24__N_1348[19]), 
          .C0(n20388), .Z(n4440)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i15 (.D(intgOut0_28__N_1629[15]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i15.GSR = "ENABLED";
    FD1P3IX intgOut3_i14 (.D(intgOut0_28__N_1629[14]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i14.GSR = "ENABLED";
    FD1P3IX intgOut3_i13 (.D(intgOut0_28__N_1629[13]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i13.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i19 (.BLUT(subIn2_24__N_1535[18]), .ALUT(subIn2_24__N_1348[18]), 
          .C0(n20388), .Z(n4441)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i12 (.D(intgOut0_28__N_1629[12]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i12.GSR = "ENABLED";
    FD1P3IX intgOut3_i11 (.D(intgOut0_28__N_1629[11]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i11.GSR = "ENABLED";
    FD1P3IX intgOut3_i10 (.D(intgOut0_28__N_1629[10]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i10.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i18 (.BLUT(subIn2_24__N_1535[17]), .ALUT(subIn2_24__N_1348[17]), 
          .C0(n20388), .Z(n4442)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i9 (.D(intgOut0_28__N_1629[9]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i9.GSR = "ENABLED";
    FD1P3IX intgOut3_i8 (.D(intgOut0_28__N_1629[8]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i8.GSR = "ENABLED";
    FD1P3IX intgOut3_i7 (.D(intgOut0_28__N_1629[7]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i7.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i17 (.BLUT(subIn2_24__N_1535[16]), .ALUT(subIn2_24__N_1348[16]), 
          .C0(n20388), .Z(n4443)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i6 (.D(intgOut0_28__N_1629[6]), .SP(clk_N_875_enable_303), 
            .CD(n14388), .CK(clk_N_875), .Q(intgOut3[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i6.GSR = "ENABLED";
    FD1P3IX intgOut3_i5 (.D(addOut[5]), .SP(clk_N_875_enable_303), .CD(n14382), 
            .CK(clk_N_875), .Q(intgOut3[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i5.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i16 (.BLUT(subIn2_24__N_1535[15]), .ALUT(subIn2_24__N_1348[15]), 
          .C0(n20388), .Z(n4444)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut3_i4 (.D(addOut[4]), .SP(clk_N_875_enable_303), .CD(n14382), 
            .CK(clk_N_875), .Q(intgOut3[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i4.GSR = "ENABLED";
    FD1P3IX intgOut3_i3 (.D(addOut[3]), .SP(clk_N_875_enable_303), .CD(n14382), 
            .CK(clk_N_875), .Q(intgOut3[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i3.GSR = "ENABLED";
    FD1P3IX intgOut3_i2 (.D(addOut[2]), .SP(clk_N_875_enable_303), .CD(n14382), 
            .CK(clk_N_875), .Q(intgOut3[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i2.GSR = "ENABLED";
    FD1P3IX intgOut3_i1 (.D(addOut[1]), .SP(clk_N_875_enable_303), .CD(n14382), 
            .CK(clk_N_875), .Q(intgOut3[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut3_i1.GSR = "ENABLED";
    FD1P3IX intgOut2_i28 (.D(intgOut0_28__N_1629[28]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i28.GSR = "ENABLED";
    CCU2D add_15129_6 (.A0(speed_set_m4[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18295), .COUT(n18296));
    defparam add_15129_6.INIT0 = 16'h5aaa;
    defparam add_15129_6.INIT1 = 16'h5aaa;
    defparam add_15129_6.INJECT1_0 = "NO";
    defparam add_15129_6.INJECT1_1 = "NO";
    PFUMX subIn2_24__I_0_rep_1_i15 (.BLUT(subIn2_24__N_1535[14]), .ALUT(subIn2_24__N_1348[14]), 
          .C0(n20388), .Z(n4445)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i27 (.D(intgOut0_28__N_1629[27]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i27.GSR = "ENABLED";
    FD1P3IX intgOut2_i26 (.D(intgOut0_28__N_1629[26]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i26.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i14 (.BLUT(subIn2_24__N_1535[13]), .ALUT(subIn2_24__N_1348[13]), 
          .C0(n20388), .Z(n4446)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i25 (.D(intgOut0_28__N_1629[25]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i25.GSR = "ENABLED";
    FD1P3IX intgOut2_i24 (.D(intgOut0_28__N_1629[24]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i24.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i12 (.BLUT(subIn2_24__N_1535[11]), .ALUT(subIn2_24__N_1348[11]), 
          .C0(n20388), .Z(n4448)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX subIn2_24__I_0_rep_1_i11 (.BLUT(subIn2_24__N_1535[10]), .ALUT(subIn2_24__N_1348[10]), 
          .C0(n20388), .Z(n4449)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX subIn2_24__I_0_rep_1_i7 (.BLUT(subIn2_24__N_1535[6]), .ALUT(subIn2_24__N_1348[6]), 
          .C0(n20388), .Z(n4453)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i23 (.D(intgOut0_28__N_1629[23]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i23.GSR = "ENABLED";
    FD1P3IX intgOut2_i22 (.D(intgOut0_28__N_1629[22]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i22.GSR = "ENABLED";
    FD1P3IX intgOut2_i21 (.D(intgOut0_28__N_1629[21]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i21.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i6 (.BLUT(subIn2_24__N_1535[5]), .ALUT(subIn2_24__N_1348[5]), 
          .C0(n20388), .Z(n4454)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX subIn2_24__I_0_rep_1_i5 (.BLUT(subIn2_24__N_1535[4]), .ALUT(subIn2_24__N_1348[4]), 
          .C0(n20388), .Z(n4455)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i20 (.D(intgOut0_28__N_1629[20]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i20.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i3 (.BLUT(subIn2_24__N_1535[2]), .ALUT(subIn2_24__N_1348[2]), 
          .C0(n20388), .Z(n4457)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX subIn2_24__I_0_rep_1_i2 (.BLUT(subIn2_24__N_1535[1]), .ALUT(subIn2_24__N_1348[1]), 
          .C0(n20388), .Z(n4458)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i19 (.D(intgOut0_28__N_1629[19]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i19.GSR = "ENABLED";
    FD1P3IX intgOut2_i18 (.D(intgOut0_28__N_1629[18]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i18.GSR = "ENABLED";
    FD1P3IX intgOut2_i17 (.D(intgOut0_28__N_1629[17]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i17.GSR = "ENABLED";
    PFUMX subIn2_24__I_0_rep_1_i1 (.BLUT(subIn2_24__N_1535[0]), .ALUT(subIn2_24__N_1348[0]), 
          .C0(n20388), .Z(n4459)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i22 (.BLUT(n558[21]), .ALUT(n678[21]), .C0(n20157), 
          .Z(addIn2_28__N_1571[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i16 (.D(intgOut0_28__N_1629[16]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i16.GSR = "ENABLED";
    FD1P3IX intgOut2_i15 (.D(intgOut0_28__N_1629[15]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i15.GSR = "ENABLED";
    FD1P3IX intgOut2_i14 (.D(intgOut0_28__N_1629[14]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i14.GSR = "ENABLED";
    FD1P3IX intgOut2_i13 (.D(intgOut0_28__N_1629[13]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i13.GSR = "ENABLED";
    PFUMX mux_140_i23 (.BLUT(n558[22]), .ALUT(n678[22]), .C0(n20157), 
          .Z(addIn2_28__N_1571[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i12 (.D(intgOut0_28__N_1629[12]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i12.GSR = "ENABLED";
    PFUMX mux_140_i2 (.BLUT(n558[1]), .ALUT(n678[1]), .C0(n20157), .Z(addIn2_28__N_1571[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i11 (.D(intgOut0_28__N_1629[11]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i11.GSR = "ENABLED";
    FD1P3IX intgOut2_i10 (.D(intgOut0_28__N_1629[10]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i10.GSR = "ENABLED";
    FD1P3IX intgOut2_i9 (.D(intgOut0_28__N_1629[9]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i9.GSR = "ENABLED";
    PFUMX mux_140_i24 (.BLUT(n558[23]), .ALUT(n678[23]), .C0(n20157), 
          .Z(addIn2_28__N_1571[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i8 (.D(intgOut0_28__N_1629[8]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i8.GSR = "ENABLED";
    CCU2D add_15129_4 (.A0(speed_set_m4[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18294), .COUT(n18295));
    defparam add_15129_4.INIT0 = 16'h5555;
    defparam add_15129_4.INIT1 = 16'h5aaa;
    defparam add_15129_4.INJECT1_0 = "NO";
    defparam add_15129_4.INJECT1_1 = "NO";
    FD1P3IX intgOut2_i7 (.D(intgOut0_28__N_1629[7]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i7.GSR = "ENABLED";
    PFUMX mux_140_i3 (.BLUT(n558[2]), .ALUT(n678[2]), .C0(n20157), .Z(addIn2_28__N_1571[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i6 (.D(intgOut0_28__N_1629[6]), .SP(clk_N_875_enable_392), 
            .CD(n14360), .CK(clk_N_875), .Q(intgOut2[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i6.GSR = "ENABLED";
    FD1P3IX intgOut2_i5 (.D(addOut[5]), .SP(clk_N_875_enable_392), .CD(n15143), 
            .CK(clk_N_875), .Q(intgOut2[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i5.GSR = "ENABLED";
    PFUMX mux_140_i25 (.BLUT(n558[24]), .ALUT(n678[24]), .C0(n20157), 
          .Z(addIn2_28__N_1571[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i4 (.BLUT(n558[3]), .ALUT(n678[3]), .C0(n20157), .Z(addIn2_28__N_1571[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i4 (.D(addOut[4]), .SP(clk_N_875_enable_392), .CD(n15143), 
            .CK(clk_N_875), .Q(intgOut2[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i4.GSR = "ENABLED";
    FD1P3IX intgOut2_i3 (.D(addOut[3]), .SP(clk_N_875_enable_392), .CD(n15143), 
            .CK(clk_N_875), .Q(intgOut2[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i3.GSR = "ENABLED";
    CCU2D add_15129_2 (.A0(speed_set_m4[1]), .B0(speed_set_m4[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18294));
    defparam add_15129_2.INIT0 = 16'h1000;
    defparam add_15129_2.INIT1 = 16'h5555;
    defparam add_15129_2.INJECT1_0 = "NO";
    defparam add_15129_2.INJECT1_1 = "NO";
    PFUMX mux_140_i26 (.BLUT(n558[25]), .ALUT(n678[25]), .C0(n20157), 
          .Z(addIn2_28__N_1571[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i2 (.D(addOut[2]), .SP(clk_N_875_enable_392), .CD(n15143), 
            .CK(clk_N_875), .Q(intgOut2[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i2.GSR = "ENABLED";
    FD1P3IX intgOut2_i1 (.D(addOut[1]), .SP(clk_N_875_enable_392), .CD(n15143), 
            .CK(clk_N_875), .Q(intgOut2[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i1.GSR = "ENABLED";
    PFUMX mux_140_i5 (.BLUT(n558[4]), .ALUT(n678[4]), .C0(n20157), .Z(addIn2_28__N_1571[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut1_i28 (.D(intgOut0_28__N_1629[28]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i28.GSR = "ENABLED";
    FD1P3IX intgOut1_i27 (.D(intgOut0_28__N_1629[27]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i27.GSR = "ENABLED";
    PFUMX mux_140_i27 (.BLUT(n558[26]), .ALUT(n678[26]), .C0(n20157), 
          .Z(addIn2_28__N_1571[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i13716_3_lut_4_lut (.A(n21465), .B(n21466), .C(n4_adj_2356), 
         .D(n3632), .Z(n16301)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i13716_3_lut_4_lut.init = 16'hfeee;
    FD1P3IX intgOut1_i26 (.D(intgOut0_28__N_1629[26]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i26.GSR = "ENABLED";
    FD1P3IX intgOut1_i25 (.D(intgOut0_28__N_1629[25]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i25.GSR = "ENABLED";
    FD1P3IX intgOut1_i24 (.D(intgOut0_28__N_1629[24]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i24.GSR = "ENABLED";
    FD1P3IX intgOut1_i23 (.D(intgOut0_28__N_1629[23]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i23.GSR = "ENABLED";
    FD1P3IX intgOut1_i22 (.D(intgOut0_28__N_1629[22]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i22.GSR = "ENABLED";
    FD1P3IX intgOut1_i21 (.D(intgOut0_28__N_1629[21]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i21.GSR = "ENABLED";
    FD1P3IX intgOut1_i20 (.D(intgOut0_28__N_1629[20]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i20.GSR = "ENABLED";
    FD1P3IX intgOut1_i19 (.D(intgOut0_28__N_1629[19]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i19.GSR = "ENABLED";
    LUT4 i1_3_lut_adj_137 (.A(n1343[15]), .B(n2305[6]), .C(n9_adj_2373), 
         .Z(n1502[6])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_137.init = 16'h8a8a;
    FD1P3IX intgOut1_i18 (.D(intgOut0_28__N_1629[18]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i18.GSR = "ENABLED";
    FD1P3IX intgOut1_i17 (.D(intgOut0_28__N_1629[17]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i17.GSR = "ENABLED";
    FD1P3IX intgOut1_i16 (.D(intgOut0_28__N_1629[16]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i16.GSR = "ENABLED";
    FD1P3IX intgOut1_i15 (.D(intgOut0_28__N_1629[15]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i15.GSR = "ENABLED";
    FD1P3IX intgOut1_i14 (.D(intgOut0_28__N_1629[14]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i14.GSR = "ENABLED";
    FD1P3IX intgOut1_i13 (.D(intgOut0_28__N_1629[13]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i13.GSR = "ENABLED";
    FD1P3IX intgOut1_i12 (.D(intgOut0_28__N_1629[12]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i12.GSR = "ENABLED";
    PFUMX mux_140_i6 (.BLUT(n558[5]), .ALUT(n678[5]), .C0(n20157), .Z(addIn2_28__N_1571[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut1_i11 (.D(intgOut0_28__N_1629[11]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i11.GSR = "ENABLED";
    PFUMX mux_140_i7 (.BLUT(n558[6]), .ALUT(n678[6]), .C0(n20157), .Z(addIn2_28__N_1571[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut1_i10 (.D(intgOut0_28__N_1629[10]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i10.GSR = "ENABLED";
    FD1P3IX intgOut1_i9 (.D(intgOut0_28__N_1629[9]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i9.GSR = "ENABLED";
    FD1P3IX intgOut1_i8 (.D(intgOut0_28__N_1629[8]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i8.GSR = "ENABLED";
    FD1P3IX intgOut1_i7 (.D(intgOut0_28__N_1629[7]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i7.GSR = "ENABLED";
    CCU2D add_15133_15 (.A0(speed_set_m4[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18486), .COUT(n18487));
    defparam add_15133_15.INIT0 = 16'hf555;
    defparam add_15133_15.INIT1 = 16'hf555;
    defparam add_15133_15.INJECT1_0 = "NO";
    defparam add_15133_15.INJECT1_1 = "NO";
    CCU2D add_15133_13 (.A0(speed_set_m4[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18485), .COUT(n18486));
    defparam add_15133_13.INIT0 = 16'hf555;
    defparam add_15133_13.INIT1 = 16'hf555;
    defparam add_15133_13.INJECT1_0 = "NO";
    defparam add_15133_13.INJECT1_1 = "NO";
    FD1P3IX intgOut1_i6 (.D(intgOut0_28__N_1629[6]), .SP(clk_N_875_enable_359), 
            .CD(n14332), .CK(clk_N_875), .Q(intgOut1[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i6.GSR = "ENABLED";
    FD1P3IX intgOut1_i5 (.D(addOut[5]), .SP(clk_N_875_enable_359), .CD(n15130), 
            .CK(clk_N_875), .Q(intgOut1[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i5.GSR = "ENABLED";
    CCU2D add_15133_11 (.A0(speed_set_m4[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18484), .COUT(n18485));
    defparam add_15133_11.INIT0 = 16'hf555;
    defparam add_15133_11.INIT1 = 16'hf555;
    defparam add_15133_11.INJECT1_0 = "NO";
    defparam add_15133_11.INJECT1_1 = "NO";
    FD1P3IX intgOut1_i4 (.D(addOut[4]), .SP(clk_N_875_enable_359), .CD(n15130), 
            .CK(clk_N_875), .Q(intgOut1[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i4.GSR = "ENABLED";
    FD1P3IX intgOut1_i3 (.D(addOut[3]), .SP(clk_N_875_enable_359), .CD(n15130), 
            .CK(clk_N_875), .Q(intgOut1[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i3.GSR = "ENABLED";
    FD1P3IX intgOut1_i2 (.D(addOut[2]), .SP(clk_N_875_enable_359), .CD(n15130), 
            .CK(clk_N_875), .Q(intgOut1[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i2.GSR = "ENABLED";
    FD1P3IX intgOut1_i1 (.D(addOut[1]), .SP(clk_N_875_enable_359), .CD(n15130), 
            .CK(clk_N_875), .Q(intgOut1[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut1_i1.GSR = "ENABLED";
    FD1P3IX intgOut0_i28 (.D(intgOut0_28__N_1629[28]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i28.GSR = "ENABLED";
    FD1P3IX intgOut0_i27 (.D(intgOut0_28__N_1629[27]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i27.GSR = "ENABLED";
    FD1P3IX intgOut0_i26 (.D(intgOut0_28__N_1629[26]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i26.GSR = "ENABLED";
    FD1P3IX intgOut0_i25 (.D(intgOut0_28__N_1629[25]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i25.GSR = "ENABLED";
    FD1P3IX intgOut0_i24 (.D(intgOut0_28__N_1629[24]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i24.GSR = "ENABLED";
    FD1P3IX intgOut0_i23 (.D(intgOut0_28__N_1629[23]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i23.GSR = "ENABLED";
    FD1P3IX intgOut0_i22 (.D(intgOut0_28__N_1629[22]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i22.GSR = "ENABLED";
    FD1P3IX intgOut0_i21 (.D(intgOut0_28__N_1629[21]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i21.GSR = "ENABLED";
    FD1P3IX intgOut0_i20 (.D(intgOut0_28__N_1629[20]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i20.GSR = "ENABLED";
    FD1P3IX intgOut0_i19 (.D(intgOut0_28__N_1629[19]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i19.GSR = "ENABLED";
    FD1P3IX intgOut0_i18 (.D(intgOut0_28__N_1629[18]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i18.GSR = "ENABLED";
    FD1P3IX intgOut0_i17 (.D(intgOut0_28__N_1629[17]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i17.GSR = "ENABLED";
    PFUMX mux_140_i28 (.BLUT(n558[27]), .ALUT(n678[27]), .C0(n20157), 
          .Z(addIn2_28__N_1571[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut0_i16 (.D(intgOut0_28__N_1629[16]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i16.GSR = "ENABLED";
    FD1P3IX intgOut0_i15 (.D(intgOut0_28__N_1629[15]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i15.GSR = "ENABLED";
    FD1P3IX intgOut0_i14 (.D(intgOut0_28__N_1629[14]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i14.GSR = "ENABLED";
    CCU2D add_211_3 (.A0(Out0[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18242), 
          .COUT(n18243), .S0(n1301[1]), .S1(n1301[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_3.INIT0 = 16'h5aaa;
    defparam add_211_3.INIT1 = 16'h5aaa;
    defparam add_211_3.INJECT1_0 = "NO";
    defparam add_211_3.INJECT1_1 = "NO";
    FD1P3IX intgOut0_i13 (.D(intgOut0_28__N_1629[13]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i13.GSR = "ENABLED";
    FD1P3IX intgOut0_i12 (.D(intgOut0_28__N_1629[12]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i12.GSR = "ENABLED";
    FD1P3IX intgOut0_i11 (.D(intgOut0_28__N_1629[11]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i11.GSR = "ENABLED";
    FD1P3IX intgOut0_i10 (.D(intgOut0_28__N_1629[10]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i10.GSR = "ENABLED";
    FD1P3IX intgOut0_i9 (.D(intgOut0_28__N_1629[9]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i9.GSR = "ENABLED";
    FD1P3IX intgOut0_i8 (.D(intgOut0_28__N_1629[8]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i8.GSR = "ENABLED";
    FD1P3IX intgOut0_i7 (.D(intgOut0_28__N_1629[7]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i7.GSR = "ENABLED";
    FD1P3IX intgOut0_i6 (.D(intgOut0_28__N_1629[6]), .SP(clk_N_875_enable_387), 
            .CD(n14304), .CK(clk_N_875), .Q(intgOut0[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i6.GSR = "ENABLED";
    FD1P3IX intgOut0_i5 (.D(addOut[5]), .SP(clk_N_875_enable_387), .CD(n14299), 
            .CK(clk_N_875), .Q(intgOut0[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i5.GSR = "ENABLED";
    FD1P3IX intgOut0_i4 (.D(addOut[4]), .SP(clk_N_875_enable_387), .CD(n14299), 
            .CK(clk_N_875), .Q(intgOut0[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i4.GSR = "ENABLED";
    FD1P3IX intgOut0_i3 (.D(addOut[3]), .SP(clk_N_875_enable_387), .CD(n14299), 
            .CK(clk_N_875), .Q(intgOut0[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i3.GSR = "ENABLED";
    FD1P3IX intgOut0_i2 (.D(addOut[2]), .SP(clk_N_875_enable_387), .CD(n14299), 
            .CK(clk_N_875), .Q(intgOut0[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i2.GSR = "ENABLED";
    FD1P3IX intgOut0_i1 (.D(addOut[1]), .SP(clk_N_875_enable_387), .CD(n14299), 
            .CK(clk_N_875), .Q(intgOut0[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut0_i1.GSR = "ENABLED";
    LUT4 i2_2_lut_adj_138 (.A(n1343[5]), .B(n1343[8]), .Z(n8_adj_2383)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_138.init = 16'heeee;
    CCU2D add_15133_9 (.A0(speed_set_m4[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18483), .COUT(n18484));
    defparam add_15133_9.INIT0 = 16'hf555;
    defparam add_15133_9.INIT1 = 16'hf555;
    defparam add_15133_9.INJECT1_0 = "NO";
    defparam add_15133_9.INJECT1_1 = "NO";
    PFUMX mux_140_i8 (.BLUT(n558[7]), .ALUT(n678[7]), .C0(n20157), .Z(addIn2_28__N_1571[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_211_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Out0[13]), .B1(n18759), .C1(n18760), .D1(Out0[28]), .COUT(n18242), 
          .S1(n1301[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(334[17:21])
    defparam add_211_1.INIT0 = 16'hF000;
    defparam add_211_1.INIT1 = 16'h56aa;
    defparam add_211_1.INJECT1_0 = "NO";
    defparam add_211_1.INJECT1_1 = "NO";
    PFUMX mux_140_i29 (.BLUT(n558[28]), .ALUT(n678[28]), .C0(n20157), 
          .Z(addIn2_28__N_1571[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i9 (.BLUT(n558[8]), .ALUT(n678[8]), .C0(n20157), .Z(addIn2_28__N_1571[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i10 (.BLUT(n558[9]), .ALUT(n678[9]), .C0(n20157), .Z(addIn2_28__N_1571[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i11 (.BLUT(n558[10]), .ALUT(n678[10]), .C0(n20157), 
          .Z(addIn2_28__N_1571[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_1212_23 (.A0(n5473), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18241), 
          .S0(n2373[21]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_23.INIT0 = 16'hf555;
    defparam add_1212_23.INIT1 = 16'h0000;
    defparam add_1212_23.INJECT1_0 = "NO";
    defparam add_1212_23.INJECT1_1 = "NO";
    PFUMX mux_140_i12 (.BLUT(n558[11]), .ALUT(n678[11]), .C0(n20157), 
          .Z(addIn2_28__N_1571[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15138_21 (.A0(speed_set_m3[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18633), .S1(n49));
    defparam add_15138_21.INIT0 = 16'h5555;
    defparam add_15138_21.INIT1 = 16'h0000;
    defparam add_15138_21.INJECT1_0 = "NO";
    defparam add_15138_21.INJECT1_1 = "NO";
    PFUMX mux_140_i13 (.BLUT(n558[12]), .ALUT(n678[12]), .C0(n20157), 
          .Z(addIn2_28__N_1571[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15138_19 (.A0(speed_set_m3[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18632), .COUT(n18633));
    defparam add_15138_19.INIT0 = 16'hf555;
    defparam add_15138_19.INIT1 = 16'hf555;
    defparam add_15138_19.INJECT1_0 = "NO";
    defparam add_15138_19.INJECT1_1 = "NO";
    CCU2D add_15138_17 (.A0(speed_set_m3[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18631), .COUT(n18632));
    defparam add_15138_17.INIT0 = 16'hf555;
    defparam add_15138_17.INIT1 = 16'hf555;
    defparam add_15138_17.INJECT1_0 = "NO";
    defparam add_15138_17.INJECT1_1 = "NO";
    CCU2D add_15138_15 (.A0(speed_set_m3[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18630), .COUT(n18631));
    defparam add_15138_15.INIT0 = 16'hf555;
    defparam add_15138_15.INIT1 = 16'hf555;
    defparam add_15138_15.INJECT1_0 = "NO";
    defparam add_15138_15.INJECT1_1 = "NO";
    CCU2D add_15138_13 (.A0(speed_set_m3[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18629), .COUT(n18630));
    defparam add_15138_13.INIT0 = 16'hf555;
    defparam add_15138_13.INIT1 = 16'hf555;
    defparam add_15138_13.INJECT1_0 = "NO";
    defparam add_15138_13.INJECT1_1 = "NO";
    CCU2D add_15138_11 (.A0(speed_set_m3[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18628), .COUT(n18629));
    defparam add_15138_11.INIT0 = 16'hf555;
    defparam add_15138_11.INIT1 = 16'hf555;
    defparam add_15138_11.INJECT1_0 = "NO";
    defparam add_15138_11.INJECT1_1 = "NO";
    CCU2D add_15138_9 (.A0(speed_set_m3[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18627), .COUT(n18628));
    defparam add_15138_9.INIT0 = 16'hf555;
    defparam add_15138_9.INIT1 = 16'hf555;
    defparam add_15138_9.INJECT1_0 = "NO";
    defparam add_15138_9.INJECT1_1 = "NO";
    LUT4 mux_1222_i1_3_lut_4_lut (.A(n16496), .B(n42), .C(speed_set_m2[0]), 
         .D(speed_set_m3[0]), .Z(n5345)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(136[23] 137[50])
    defparam mux_1222_i1_3_lut_4_lut.init = 16'hfb40;
    CCU2D add_15138_7 (.A0(speed_set_m3[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18626), .COUT(n18627));
    defparam add_15138_7.INIT0 = 16'hf555;
    defparam add_15138_7.INIT1 = 16'hf555;
    defparam add_15138_7.INJECT1_0 = "NO";
    defparam add_15138_7.INJECT1_1 = "NO";
    PFUMX mux_140_i14 (.BLUT(n558[13]), .ALUT(n678[13]), .C0(n20157), 
          .Z(addIn2_28__N_1571[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i15 (.BLUT(n558[14]), .ALUT(n678[14]), .C0(n20157), 
          .Z(addIn2_28__N_1571[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15138_5 (.A0(speed_set_m3[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18625), .COUT(n18626));
    defparam add_15138_5.INIT0 = 16'hf555;
    defparam add_15138_5.INIT1 = 16'hf555;
    defparam add_15138_5.INJECT1_0 = "NO";
    defparam add_15138_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_139 (.A(n1343[3]), .B(n1343[2]), .C(n1343[1]), .D(n1343[0]), 
         .Z(n4_adj_2384)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_139.init = 16'haaa8;
    CCU2D add_15133_7 (.A0(speed_set_m4[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18482), .COUT(n18483));
    defparam add_15133_7.INIT0 = 16'hf555;
    defparam add_15133_7.INIT1 = 16'hf555;
    defparam add_15133_7.INJECT1_0 = "NO";
    defparam add_15133_7.INJECT1_1 = "NO";
    CCU2D add_15133_5 (.A0(speed_set_m4[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18481), .COUT(n18482));
    defparam add_15133_5.INIT0 = 16'hf555;
    defparam add_15133_5.INIT1 = 16'hf555;
    defparam add_15133_5.INJECT1_0 = "NO";
    defparam add_15133_5.INJECT1_1 = "NO";
    CCU2D add_15133_3 (.A0(speed_set_m4[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m4[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18480), .COUT(n18481));
    defparam add_15133_3.INIT0 = 16'hf555;
    defparam add_15133_3.INIT1 = 16'hf555;
    defparam add_15133_3.INJECT1_0 = "NO";
    defparam add_15133_3.INJECT1_1 = "NO";
    CCU2D add_15138_3 (.A0(speed_set_m3[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18624), .COUT(n18625));
    defparam add_15138_3.INIT0 = 16'hf555;
    defparam add_15138_3.INIT1 = 16'hf555;
    defparam add_15138_3.INJECT1_0 = "NO";
    defparam add_15138_3.INJECT1_1 = "NO";
    CCU2D add_15133_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m4[0]), .B1(speed_set_m4[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18480));
    defparam add_15133_1.INIT0 = 16'hF000;
    defparam add_15133_1.INIT1 = 16'ha666;
    defparam add_15133_1.INJECT1_0 = "NO";
    defparam add_15133_1.INJECT1_1 = "NO";
    CCU2D add_15138_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m3[0]), .B1(speed_set_m3[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18624));
    defparam add_15138_1.INIT0 = 16'hF000;
    defparam add_15138_1.INIT1 = 16'ha666;
    defparam add_15138_1.INJECT1_0 = "NO";
    defparam add_15138_1.INJECT1_1 = "NO";
    LUT4 i14060_3_lut_4_lut (.A(n21465), .B(n21466), .C(n4_adj_2341), 
         .D(n3728), .Z(n16670)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(234[73:80])
    defparam i14060_3_lut_4_lut.init = 16'hfeee;
    CCU2D addOut_2126_add_4_29 (.A0(multOut[27]), .B0(n16420), .C0(addOut[27]), 
          .D0(addIn2_28__N_1441[27]), .A1(multOut[28]), .B1(n16420), .C1(addOut[28]), 
          .D1(addIn2_28__N_1441[28]), .CIN(n18420), .S0(n121[27]), .S1(n121[28]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_29.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_29.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_29.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_29.INJECT1_1 = "NO";
    PFUMX mux_140_i16 (.BLUT(n558[15]), .ALUT(n678[15]), .C0(n20157), 
          .Z(addIn2_28__N_1571[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D addOut_2126_add_4_27 (.A0(multOut[25]), .B0(n16420), .C0(addOut[25]), 
          .D0(addIn2_28__N_1441[25]), .A1(multOut[26]), .B1(n16420), .C1(addOut[26]), 
          .D1(addIn2_28__N_1441[26]), .CIN(n18419), .COUT(n18420), .S0(n121[25]), 
          .S1(n121[26]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_27.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_27.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_27.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_27.INJECT1_1 = "NO";
    LUT4 i17233_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut_4_lut (.A(n21499), .B(ss[0]), 
         .C(ss[2]), .D(ss[1]), .Z(n20374)) /* synthesis lut_function=(!(A+(B (C (D))+!B !(C+(D))))) */ ;
    defparam i17233_2_lut_3_lut_4_lut_2_lut_3_lut_4_lut_4_lut.init = 16'h1554;
    CCU2D add_1212_21 (.A0(n5471), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5473), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18240), 
          .COUT(n18241), .S0(n2373[19]), .S1(n2373[20]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_21.INIT0 = 16'hf555;
    defparam add_1212_21.INIT1 = 16'hf555;
    defparam add_1212_21.INJECT1_0 = "NO";
    defparam add_1212_21.INJECT1_1 = "NO";
    PFUMX mux_140_i17 (.BLUT(n558[16]), .ALUT(n678[16]), .C0(n20157), 
          .Z(addIn2_28__N_1571[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i18 (.BLUT(n558[17]), .ALUT(n678[17]), .C0(n20157), 
          .Z(addIn2_28__N_1571[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_1212_19 (.A0(n5467), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5469), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18239), 
          .COUT(n18240), .S0(n2373[17]), .S1(n2373[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_19.INIT0 = 16'hf555;
    defparam add_1212_19.INIT1 = 16'hf555;
    defparam add_1212_19.INJECT1_0 = "NO";
    defparam add_1212_19.INJECT1_1 = "NO";
    PFUMX mux_140_i19 (.BLUT(n558[18]), .ALUT(n678[18]), .C0(n20157), 
          .Z(addIn2_28__N_1571[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15130_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18613), 
          .S0(n3728));
    defparam add_15130_cout.INIT0 = 16'h0000;
    defparam add_15130_cout.INIT1 = 16'h0000;
    defparam add_15130_cout.INJECT1_0 = "NO";
    defparam add_15130_cout.INJECT1_1 = "NO";
    PFUMX mux_140_i20 (.BLUT(n558[19]), .ALUT(n678[19]), .C0(n20157), 
          .Z(addIn2_28__N_1571[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_140_i21 (.BLUT(n558[20]), .ALUT(n678[20]), .C0(n20157), 
          .Z(addIn2_28__N_1571[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15130_20 (.A0(speed_set_m3[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18612), .COUT(n18613));
    defparam add_15130_20.INIT0 = 16'h5aaa;
    defparam add_15130_20.INIT1 = 16'h0aaa;
    defparam add_15130_20.INJECT1_0 = "NO";
    defparam add_15130_20.INJECT1_1 = "NO";
    CCU2D add_15130_18 (.A0(speed_set_m3[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18611), .COUT(n18612));
    defparam add_15130_18.INIT0 = 16'h5aaa;
    defparam add_15130_18.INIT1 = 16'h5aaa;
    defparam add_15130_18.INJECT1_0 = "NO";
    defparam add_15130_18.INJECT1_1 = "NO";
    CCU2D add_15130_16 (.A0(speed_set_m3[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18610), .COUT(n18611));
    defparam add_15130_16.INIT0 = 16'h5aaa;
    defparam add_15130_16.INIT1 = 16'h5aaa;
    defparam add_15130_16.INJECT1_0 = "NO";
    defparam add_15130_16.INJECT1_1 = "NO";
    PFUMX mux_140_i1 (.BLUT(n558[0]), .ALUT(n678[0]), .C0(n20157), .Z(addIn2_28__N_1571[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15130_14 (.A0(speed_set_m3[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18609), .COUT(n18610));
    defparam add_15130_14.INIT0 = 16'h5555;
    defparam add_15130_14.INIT1 = 16'h5aaa;
    defparam add_15130_14.INJECT1_0 = "NO";
    defparam add_15130_14.INJECT1_1 = "NO";
    CCU2D add_15130_12 (.A0(speed_set_m3[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18608), .COUT(n18609));
    defparam add_15130_12.INIT0 = 16'h5aaa;
    defparam add_15130_12.INIT1 = 16'h5aaa;
    defparam add_15130_12.INJECT1_0 = "NO";
    defparam add_15130_12.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_347_3_lut_4_lut (.A(ss[0]), .B(ss[1]), .C(ss[2]), 
         .D(n21499), .Z(n21448)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_2_lut_rep_347_3_lut_4_lut.init = 16'h0060;
    LUT4 i1_3_lut_adj_140 (.A(n1343[15]), .B(n2305[5]), .C(n9_adj_2373), 
         .Z(n1502[5])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_140.init = 16'h8a8a;
    PFUMX mux_137_i22 (.BLUT(n588[21]), .ALUT(intgOut3[21]), .C0(n21420), 
          .Z(n618[21])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_15130_10 (.A0(speed_set_m3[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18607), .COUT(n18608));
    defparam add_15130_10.INIT0 = 16'h5555;
    defparam add_15130_10.INIT1 = 16'h5555;
    defparam add_15130_10.INJECT1_0 = "NO";
    defparam add_15130_10.INJECT1_1 = "NO";
    CCU2D add_15130_8 (.A0(speed_set_m3[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18606), .COUT(n18607));
    defparam add_15130_8.INIT0 = 16'h5aaa;
    defparam add_15130_8.INIT1 = 16'h5555;
    defparam add_15130_8.INJECT1_0 = "NO";
    defparam add_15130_8.INJECT1_1 = "NO";
    CCU2D add_15130_6 (.A0(speed_set_m3[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18605), .COUT(n18606));
    defparam add_15130_6.INIT0 = 16'h5aaa;
    defparam add_15130_6.INIT1 = 16'h5aaa;
    defparam add_15130_6.INJECT1_0 = "NO";
    defparam add_15130_6.INJECT1_1 = "NO";
    CCU2D add_15130_4 (.A0(speed_set_m3[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18604), .COUT(n18605));
    defparam add_15130_4.INIT0 = 16'h5555;
    defparam add_15130_4.INIT1 = 16'h5aaa;
    defparam add_15130_4.INJECT1_0 = "NO";
    defparam add_15130_4.INJECT1_1 = "NO";
    CCU2D add_1212_17 (.A0(n5463), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5465), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18238), 
          .COUT(n18239), .S0(n2373[15]), .S1(n2373[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_17.INIT0 = 16'hf555;
    defparam add_1212_17.INIT1 = 16'hf555;
    defparam add_1212_17.INJECT1_0 = "NO";
    defparam add_1212_17.INJECT1_1 = "NO";
    CCU2D add_15130_2 (.A0(speed_set_m3[1]), .B0(speed_set_m3[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m3[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18604));
    defparam add_15130_2.INIT0 = 16'h1000;
    defparam add_15130_2.INIT1 = 16'h5555;
    defparam add_15130_2.INJECT1_0 = "NO";
    defparam add_15130_2.INJECT1_1 = "NO";
    LUT4 ss_0__bdd_4_lut (.A(ss[0]), .B(ss[2]), .C(n22216), .D(ss[3]), 
         .Z(n16420)) /* synthesis lut_function=(A+(B (C+(D))+!B (C+!(D)))) */ ;
    defparam ss_0__bdd_4_lut.init = 16'hfefb;
    PFUMX mux_137_i23 (.BLUT(n588[22]), .ALUT(intgOut3[22]), .C0(n21420), 
          .Z(n618[22])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i11824_4_lut (.A(clk_N_875_enable_391), .B(n1343[15]), .C(n9_adj_2373), 
         .D(n21463), .Z(n14428)) /* synthesis lut_function=(A (((D)+!C)+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i11824_4_lut.init = 16'haa2a;
    LUT4 i1_3_lut_adj_141 (.A(n1343[15]), .B(n2305[3]), .C(n9_adj_2373), 
         .Z(n1502[3])) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_141.init = 16'h8a8a;
    PFUMX mux_137_i24 (.BLUT(n588[23]), .ALUT(intgOut3[23]), .C0(n21420), 
          .Z(n618[23])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i25 (.BLUT(n588[24]), .ALUT(intgOut3[24]), .C0(n21420), 
          .Z(n618[24])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i26 (.BLUT(n588[25]), .ALUT(intgOut3[25]), .C0(n21420), 
          .Z(n618[25])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m4_i0_i0 (.D(n2317[0]), .SP(clk_N_875_enable_391), .CD(n14437), 
            .CK(clk_N_875), .Q(PWMdut_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m4_i0_i0.GSR = "DISABLED";
    FD1P3IX dutyout_m3_i0_i0 (.D(n2305[0]), .SP(clk_N_875_enable_391), .CD(n14428), 
            .CK(clk_N_875), .Q(PWMdut_m3[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m3_i0_i0.GSR = "DISABLED";
    FD1P3IX dutyout_m2_i0_i0 (.D(n2293[0]), .SP(clk_N_875_enable_391), .CD(n14419), 
            .CK(clk_N_875), .Q(PWMdut_m2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m2_i0_i0.GSR = "DISABLED";
    PFUMX mux_137_i27 (.BLUT(n588[26]), .ALUT(intgOut3[26]), .C0(n21420), 
          .Z(n618[26])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i28 (.BLUT(n588[27]), .ALUT(intgOut3[27]), .C0(n21420), 
          .Z(n618[27])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX dutyout_m1_i0_i0 (.D(n2281[0]), .SP(clk_N_875_enable_391), .CD(n14410), 
            .CK(clk_N_875), .Q(PWMdut_m1[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam dutyout_m1_i0_i0.GSR = "DISABLED";
    CCU2D sub_16_rep_4_add_2_23 (.A0(n8_adj_2372), .B0(n16542), .C0(n5909), 
          .D0(n16223), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18593), .S0(n4510));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_23.INIT0 = 16'h0f8f;
    defparam sub_16_rep_4_add_2_23.INIT1 = 16'h0000;
    defparam sub_16_rep_4_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_21 (.A0(n4440), .B0(n11585), .C0(n5905), 
          .D0(n16223), .A1(n8_adj_2372), .B1(n16542), .C1(n5909), .D1(n16223), 
          .CIN(n18592), .COUT(n18593), .S0(n4512), .S1(n4511));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_21.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_21.INIT1 = 16'h0f8f;
    defparam sub_16_rep_4_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_21.INJECT1_1 = "NO";
    LUT4 i1827_1_lut_rep_389 (.A(ss[0]), .Z(n21490)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1827_1_lut_rep_389.init = 16'h5555;
    CCU2D sub_16_rep_4_add_2_19 (.A0(n4442), .B0(n11585), .C0(n5901), 
          .D0(n16223), .A1(n4441), .B1(n11585), .C1(n5903), .D1(n16223), 
          .CIN(n18591), .COUT(n18592), .S0(n4514), .S1(n4513));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_19.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_19.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_17 (.A0(n4444), .B0(n11585), .C0(n5897), 
          .D0(n16223), .A1(n4443), .B1(n11585), .C1(n5899), .D1(n16223), 
          .CIN(n18590), .COUT(n18591), .S0(n4516), .S1(n4515));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_17.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_17.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_17.INJECT1_1 = "NO";
    LUT4 ss_4__I_0_350_i6_2_lut_rep_364_2_lut (.A(ss[0]), .B(ss[1]), .Z(n21465)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam ss_4__I_0_350_i6_2_lut_rep_364_2_lut.init = 16'hdddd;
    CCU2D sub_16_rep_4_add_2_15 (.A0(n4446), .B0(n11585), .C0(n5893), 
          .D0(n16223), .A1(n4445), .B1(n11585), .C1(n5895), .D1(n16223), 
          .CIN(n18589), .COUT(n18590), .S0(n4518), .S1(n4517));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_15.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_15.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_13 (.A0(n4448), .B0(n11585), .C0(n5889), 
          .D0(n16223), .A1(n4447), .B1(n11585), .C1(n5891), .D1(n16223), 
          .CIN(n18588), .COUT(n18589), .S0(n4520), .S1(n4519));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_13.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_13.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_13.INJECT1_1 = "NO";
    LUT4 i17273_2_lut_rep_319_2_lut_3_lut_4_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21498), .D(ss[3]), .Z(n21420)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i17273_2_lut_rep_319_2_lut_3_lut_4_lut_4_lut.init = 16'h0200;
    PFUMX mux_137_i29 (.BLUT(n588[28]), .ALUT(intgOut3[28]), .C0(n21420), 
          .Z(n618[28])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D sub_16_rep_4_add_2_11 (.A0(n4450), .B0(n11585), .C0(n5885), 
          .D0(n16223), .A1(n4449), .B1(n11585), .C1(n5887), .D1(n16223), 
          .CIN(n18587), .COUT(n18588), .S0(n4522), .S1(n4521));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_11.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_11.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_9 (.A0(n4452), .B0(n11585), .C0(n5881), .D0(n16223), 
          .A1(n4451), .B1(n11585), .C1(n5883), .D1(n16223), .CIN(n18586), 
          .COUT(n18587), .S0(n4524), .S1(n4523));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_9.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_9.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_16_rep_4_add_2_7 (.A0(n4454), .B0(n11585), .C0(n5877), .D0(n16223), 
          .A1(n4453), .B1(n11585), .C1(n5879), .D1(n16223), .CIN(n18585), 
          .COUT(n18586), .S0(n4526), .S1(n4525));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_7.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_7.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_142 (.A(n1322[15]), .B(n2293[9]), .C(n30), .Z(n19113)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(354[4] 360[11])
    defparam i1_3_lut_adj_142.init = 16'h8a8a;
    CCU2D sub_16_rep_4_add_2_5 (.A0(n4456), .B0(n11585), .C0(n5873), .D0(n16223), 
          .A1(n4455), .B1(n11585), .C1(n5875), .D1(n16223), .CIN(n18584), 
          .COUT(n18585), .S0(n4528), .S1(n4527));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_5.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_5.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_5.INJECT1_1 = "NO";
    PFUMX mux_137_i1 (.BLUT(n588[0]), .ALUT(intgOut3[0]), .C0(n21420), 
          .Z(n618[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i5_4_lut_adj_143 (.A(n9_adj_2379), .B(n7_adj_2385), .C(n1322[10]), 
         .D(n1322[13]), .Z(n30)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut_adj_143.init = 16'h8000;
    CCU2D sub_16_rep_4_add_2_3 (.A0(n4458), .B0(n11585), .C0(n5869), .D0(n16223), 
          .A1(n4457), .B1(n11585), .C1(n5871), .D1(n16223), .CIN(n18583), 
          .COUT(n18584), .S0(n4530), .S1(n4529));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_3.INIT0 = 16'ha565;
    defparam sub_16_rep_4_add_2_3.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_3.INJECT1_1 = "NO";
    PFUMX mux_137_i2 (.BLUT(n588[1]), .ALUT(intgOut3[1]), .C0(n21420), 
          .Z(n618[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D sub_16_rep_4_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n4459), .B1(n11585), .C1(n5557), .D1(n16223), 
          .COUT(n18583), .S1(n4531));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_4_add_2_1.INIT0 = 16'h0000;
    defparam sub_16_rep_4_add_2_1.INIT1 = 16'ha565;
    defparam sub_16_rep_4_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_4_add_2_1.INJECT1_1 = "NO";
    LUT4 ss_4__I_0_358_i9_2_lut_rep_331_3_lut_4_lut_4_lut (.A(ss[0]), .B(ss[1]), 
         .C(n21494), .D(ss[3]), .Z(n21432)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam ss_4__I_0_358_i9_2_lut_rep_331_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 equal_114_i9_2_lut_rep_329_3_lut_4_lut_4_lut (.A(ss[0]), .B(ss[3]), 
         .C(n21494), .D(ss[1]), .Z(n21430)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam equal_114_i9_2_lut_rep_329_3_lut_4_lut_4_lut.init = 16'hfff7;
    PFUMX mux_137_i3 (.BLUT(n588[2]), .ALUT(intgOut3[2]), .C0(n21420), 
          .Z(n618[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1P3IX intgOut2_i0 (.D(addOut[0]), .SP(clk_N_875_enable_392), .CD(n15143), 
            .CK(clk_N_875), .Q(intgOut2[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam intgOut2_i0.GSR = "ENABLED";
    CCU2D sub_16_rep_3_add_2_23 (.A0(n2373[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18581), .S0(n4485), .S1(n4484));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_23.INIT0 = 16'h5555;
    defparam sub_16_rep_3_add_2_23.INIT1 = 16'h5555;
    defparam sub_16_rep_3_add_2_23.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_23.INJECT1_1 = "NO";
    PFUMX mux_137_i4 (.BLUT(n588[3]), .ALUT(intgOut3[3]), .C0(n21420), 
          .Z(n618[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D sub_16_rep_3_add_2_21 (.A0(n2373[19]), .B0(n4440), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18580), .COUT(n18581), .S0(n4487), .S1(n4486));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_21.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_21.INIT1 = 16'h5555;
    defparam sub_16_rep_3_add_2_21.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_21.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut (.A(ss[0]), .B(n22216), .C(n21492), .D(ss[3]), 
         .Z(multIn2[0])) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(254[3] 410[12])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0110;
    PFUMX mux_137_i5 (.BLUT(n588[4]), .ALUT(intgOut3[4]), .C0(n21420), 
          .Z(n618[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i1_2_lut_rep_390 (.A(ss[0]), .B(ss[3]), .Z(n21491)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_2_lut_rep_390.init = 16'heeee;
    LUT4 i1_2_lut_rep_337_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), 
         .D(n21494), .Z(n21438)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_2_lut_rep_337_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_144 (.A(ss[0]), .B(ss[3]), .C(ss[1]), .D(n22209), 
         .Z(n18698)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i2_3_lut_4_lut_adj_144.init = 16'h1000;
    LUT4 i1_4_lut_adj_145 (.A(n11644), .B(n19662), .C(n22216), .D(n21472), 
         .Z(clk_N_875_enable_237)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_145.init = 16'hc8c0;
    LUT4 i1_2_lut_rep_339_3_lut_4_lut (.A(ss[0]), .B(ss[3]), .C(ss[1]), 
         .D(n21494), .Z(n21440)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_2_lut_rep_339_3_lut_4_lut.init = 16'hffef;
    CCU2D sub_16_rep_3_add_2_19 (.A0(n2373[17]), .B0(n4442), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[18]), .B1(n4441), .C1(GND_net), .D1(GND_net), 
          .CIN(n18579), .COUT(n18580), .S0(n4489), .S1(n4488));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_19.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_19.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_19.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_19.INJECT1_1 = "NO";
    PFUMX mux_137_i6 (.BLUT(n588[5]), .ALUT(intgOut3[5]), .C0(n21420), 
          .Z(n618[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i7 (.BLUT(n588[6]), .ALUT(intgOut3[6]), .C0(n21420), 
          .Z(n618[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i8 (.BLUT(n588[7]), .ALUT(intgOut3[7]), .C0(n21420), 
          .Z(n618[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_146 (.A(ss[0]), .B(ss[3]), .C(ss[1]), 
         .D(n22209), .Z(n19646)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam i1_2_lut_3_lut_4_lut_adj_146.init = 16'h0100;
    PFUMX mux_137_i9 (.BLUT(n588[8]), .ALUT(intgOut3[8]), .C0(n21420), 
          .Z(n618[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    LUT4 i1_4_lut_adj_147 (.A(n1322[11]), .B(n1322[9]), .C(n10), .D(n1322[7]), 
         .Z(n7_adj_2385)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_147.init = 16'haaa8;
    FD1S3AY ss_i4_rep_410 (.D(n19674), .CK(clk_N_875), .Q(n22216));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i4_rep_410.GSR = "ENABLED";
    CCU2D sub_16_rep_3_add_2_17 (.A0(n2373[15]), .B0(n4444), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[16]), .B1(n4443), .C1(GND_net), .D1(GND_net), 
          .CIN(n18578), .COUT(n18579), .S0(n4491), .S1(n4490));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_17.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_17.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_17.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_15 (.A0(n2373[13]), .B0(n4446), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[14]), .B1(n4445), .C1(GND_net), .D1(GND_net), 
          .CIN(n18577), .COUT(n18578), .S0(n4493), .S1(n4492));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_15.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_15.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_15.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_13 (.A0(n2373[11]), .B0(n4448), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[12]), .B1(n4447), .C1(GND_net), .D1(GND_net), 
          .CIN(n18576), .COUT(n18577), .S0(n4495), .S1(n4494));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_13.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_13.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_13.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_11 (.A0(n2373[9]), .B0(n4450), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[10]), .B1(n4449), .C1(GND_net), .D1(GND_net), 
          .CIN(n18575), .COUT(n18576), .S0(n4497), .S1(n4496));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_11.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_11.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_11.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_9 (.A0(n2373[7]), .B0(n4452), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[8]), .B1(n4451), .C1(GND_net), .D1(GND_net), 
          .CIN(n18574), .COUT(n18575), .S0(n4499), .S1(n4498));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_9.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_9.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_9.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_9.INJECT1_1 = "NO";
    PFUMX mux_137_i10 (.BLUT(n588[9]), .ALUT(intgOut3[9]), .C0(n21420), 
          .Z(n618[9])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D sub_16_rep_3_add_2_7 (.A0(n2373[5]), .B0(n4454), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[6]), .B1(n4453), .C1(GND_net), .D1(GND_net), 
          .CIN(n18573), .COUT(n18574), .S0(n4501), .S1(n4500));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_7.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_7.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_7.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_5 (.A0(n2373[3]), .B0(n4456), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[4]), .B1(n4455), .C1(GND_net), .D1(GND_net), 
          .CIN(n18572), .COUT(n18573), .S0(n4503), .S1(n4502));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_5.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_5.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_5.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_3 (.A0(n2373[1]), .B0(n4458), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[2]), .B1(n4457), .C1(GND_net), .D1(GND_net), 
          .CIN(n18571), .COUT(n18572), .S0(n4505), .S1(n4504));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_3.INIT0 = 16'h5999;
    defparam sub_16_rep_3_add_2_3.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_3.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_16_rep_3_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n2373[0]), .B1(n4459), .C1(GND_net), .D1(GND_net), 
          .COUT(n18571), .S1(n4506));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(228[13:19])
    defparam sub_16_rep_3_add_2_1.INIT0 = 16'h0000;
    defparam sub_16_rep_3_add_2_1.INIT1 = 16'h5999;
    defparam sub_16_rep_3_add_2_1.INJECT1_0 = "NO";
    defparam sub_16_rep_3_add_2_1.INJECT1_1 = "NO";
    FD1S3IX ss_i2_rep_403 (.D(n14), .CK(clk_N_875), .CD(ss[4]), .Q(n22209));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(204[2] 412[9])
    defparam ss_i2_rep_403.GSR = "ENABLED";
    PFUMX mux_137_i11 (.BLUT(n588[10]), .ALUT(intgOut3[10]), .C0(n21420), 
          .Z(n618[10])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i12 (.BLUT(n588[11]), .ALUT(intgOut3[11]), .C0(n21420), 
          .Z(n618[11])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX i17353 (.BLUT(n21507), .ALUT(n21508), .C0(ss[0]), .Z(n4389));
    CCU2D add_15131_17 (.A0(speed_set_m1[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18552), .S1(n3608));
    defparam add_15131_17.INIT0 = 16'h5555;
    defparam add_15131_17.INIT1 = 16'h0000;
    defparam add_15131_17.INJECT1_0 = "NO";
    defparam add_15131_17.INJECT1_1 = "NO";
    CCU2D add_15131_15 (.A0(speed_set_m1[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18551), .COUT(n18552));
    defparam add_15131_15.INIT0 = 16'hf555;
    defparam add_15131_15.INIT1 = 16'hf555;
    defparam add_15131_15.INJECT1_0 = "NO";
    defparam add_15131_15.INJECT1_1 = "NO";
    CCU2D add_15131_13 (.A0(speed_set_m1[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18550), .COUT(n18551));
    defparam add_15131_13.INIT0 = 16'hf555;
    defparam add_15131_13.INIT1 = 16'hf555;
    defparam add_15131_13.INJECT1_0 = "NO";
    defparam add_15131_13.INJECT1_1 = "NO";
    CCU2D add_15131_11 (.A0(speed_set_m1[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18549), .COUT(n18550));
    defparam add_15131_11.INIT0 = 16'hf555;
    defparam add_15131_11.INIT1 = 16'hf555;
    defparam add_15131_11.INJECT1_0 = "NO";
    defparam add_15131_11.INJECT1_1 = "NO";
    CCU2D add_15131_9 (.A0(speed_set_m1[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18548), .COUT(n18549));
    defparam add_15131_9.INIT0 = 16'hf555;
    defparam add_15131_9.INIT1 = 16'h0aaa;
    defparam add_15131_9.INJECT1_0 = "NO";
    defparam add_15131_9.INJECT1_1 = "NO";
    CCU2D add_15131_7 (.A0(speed_set_m1[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18547), .COUT(n18548));
    defparam add_15131_7.INIT0 = 16'h0aaa;
    defparam add_15131_7.INIT1 = 16'hf555;
    defparam add_15131_7.INJECT1_0 = "NO";
    defparam add_15131_7.INJECT1_1 = "NO";
    CCU2D add_15131_5 (.A0(speed_set_m1[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18546), .COUT(n18547));
    defparam add_15131_5.INIT0 = 16'h0aaa;
    defparam add_15131_5.INIT1 = 16'h0aaa;
    defparam add_15131_5.INJECT1_0 = "NO";
    defparam add_15131_5.INJECT1_1 = "NO";
    CCU2D add_15131_3 (.A0(speed_set_m1[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m1[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18545), .COUT(n18546));
    defparam add_15131_3.INIT0 = 16'hf555;
    defparam add_15131_3.INIT1 = 16'hf555;
    defparam add_15131_3.INJECT1_0 = "NO";
    defparam add_15131_3.INJECT1_1 = "NO";
    CCU2D add_15131_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(speed_set_m1[4]), .B1(speed_set_m1[5]), .C1(GND_net), .D1(GND_net), 
          .COUT(n18545));
    defparam add_15131_1.INIT0 = 16'hF000;
    defparam add_15131_1.INIT1 = 16'ha666;
    defparam add_15131_1.INJECT1_0 = "NO";
    defparam add_15131_1.INJECT1_1 = "NO";
    CCU2D add_15132_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18544), 
          .S0(n3680));
    defparam add_15132_cout.INIT0 = 16'h0000;
    defparam add_15132_cout.INIT1 = 16'h0000;
    defparam add_15132_cout.INJECT1_0 = "NO";
    defparam add_15132_cout.INJECT1_1 = "NO";
    CCU2D add_15132_20 (.A0(speed_set_m2[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18543), .COUT(n18544));
    defparam add_15132_20.INIT0 = 16'h5aaa;
    defparam add_15132_20.INIT1 = 16'h0aaa;
    defparam add_15132_20.INJECT1_0 = "NO";
    defparam add_15132_20.INJECT1_1 = "NO";
    CCU2D add_15132_18 (.A0(speed_set_m2[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18542), .COUT(n18543));
    defparam add_15132_18.INIT0 = 16'h5aaa;
    defparam add_15132_18.INIT1 = 16'h5aaa;
    defparam add_15132_18.INJECT1_0 = "NO";
    defparam add_15132_18.INJECT1_1 = "NO";
    CCU2D add_15132_16 (.A0(speed_set_m2[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18541), .COUT(n18542));
    defparam add_15132_16.INIT0 = 16'h5aaa;
    defparam add_15132_16.INIT1 = 16'h5aaa;
    defparam add_15132_16.INJECT1_0 = "NO";
    defparam add_15132_16.INJECT1_1 = "NO";
    CCU2D add_15132_14 (.A0(speed_set_m2[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18540), .COUT(n18541));
    defparam add_15132_14.INIT0 = 16'h5555;
    defparam add_15132_14.INIT1 = 16'h5aaa;
    defparam add_15132_14.INJECT1_0 = "NO";
    defparam add_15132_14.INJECT1_1 = "NO";
    CCU2D add_15132_12 (.A0(speed_set_m2[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18539), .COUT(n18540));
    defparam add_15132_12.INIT0 = 16'h5aaa;
    defparam add_15132_12.INIT1 = 16'h5aaa;
    defparam add_15132_12.INJECT1_0 = "NO";
    defparam add_15132_12.INJECT1_1 = "NO";
    CCU2D add_15132_10 (.A0(speed_set_m2[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18538), .COUT(n18539));
    defparam add_15132_10.INIT0 = 16'h5555;
    defparam add_15132_10.INIT1 = 16'h5555;
    defparam add_15132_10.INJECT1_0 = "NO";
    defparam add_15132_10.INJECT1_1 = "NO";
    CCU2D add_15132_8 (.A0(speed_set_m2[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18537), .COUT(n18538));
    defparam add_15132_8.INIT0 = 16'h5aaa;
    defparam add_15132_8.INIT1 = 16'h5555;
    defparam add_15132_8.INJECT1_0 = "NO";
    defparam add_15132_8.INJECT1_1 = "NO";
    CCU2D add_15132_6 (.A0(speed_set_m2[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18536), .COUT(n18537));
    defparam add_15132_6.INIT0 = 16'h5aaa;
    defparam add_15132_6.INIT1 = 16'h5aaa;
    defparam add_15132_6.INJECT1_0 = "NO";
    defparam add_15132_6.INJECT1_1 = "NO";
    CCU2D add_15132_4 (.A0(speed_set_m2[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n18535), .COUT(n18536));
    defparam add_15132_4.INIT0 = 16'h5555;
    defparam add_15132_4.INIT1 = 16'h5aaa;
    defparam add_15132_4.INJECT1_0 = "NO";
    defparam add_15132_4.INJECT1_1 = "NO";
    CCU2D add_15132_2 (.A0(speed_set_m2[1]), .B0(speed_set_m2[0]), .C0(GND_net), 
          .D0(GND_net), .A1(speed_set_m2[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n18535));
    defparam add_15132_2.INIT0 = 16'h1000;
    defparam add_15132_2.INIT1 = 16'h5555;
    defparam add_15132_2.INJECT1_0 = "NO";
    defparam add_15132_2.INJECT1_1 = "NO";
    CCU2D add_1212_15 (.A0(n5459), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5461), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18237), 
          .COUT(n18238), .S0(n2373[13]), .S1(n2373[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_15.INIT0 = 16'hf555;
    defparam add_1212_15.INIT1 = 16'hf555;
    defparam add_1212_15.INJECT1_0 = "NO";
    defparam add_1212_15.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_25 (.A0(multOut[23]), .B0(n16420), .C0(addOut[23]), 
          .D0(addIn2_28__N_1441[23]), .A1(multOut[24]), .B1(n16420), .C1(addOut[24]), 
          .D1(addIn2_28__N_1441[24]), .CIN(n18418), .COUT(n18419), .S0(n121[23]), 
          .S1(n121[24]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_25.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_25.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_25.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_25.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_23 (.A0(multOut[21]), .B0(n16420), .C0(addOut[21]), 
          .D0(addIn2_28__N_1441[21]), .A1(multOut[22]), .B1(n16420), .C1(addOut[22]), 
          .D1(addIn2_28__N_1441[22]), .CIN(n18417), .COUT(n18418), .S0(n121[21]), 
          .S1(n121[22]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_23.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_23.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_23.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_23.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_21 (.A0(multOut[19]), .B0(n16420), .C0(addOut[19]), 
          .D0(addIn2_28__N_1441[19]), .A1(multOut[20]), .B1(n16420), .C1(addOut[20]), 
          .D1(addIn2_28__N_1441[20]), .CIN(n18416), .COUT(n18417), .S0(n121[19]), 
          .S1(n121[20]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_21.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_21.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_21.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_21.INJECT1_1 = "NO";
    CCU2D add_1212_13 (.A0(n5455), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5457), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18236), 
          .COUT(n18237), .S0(n2373[11]), .S1(n2373[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_13.INIT0 = 16'hf555;
    defparam add_1212_13.INIT1 = 16'hf555;
    defparam add_1212_13.INJECT1_0 = "NO";
    defparam add_1212_13.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_19 (.A0(multOut[17]), .B0(n16420), .C0(addOut[17]), 
          .D0(addIn2_28__N_1441[17]), .A1(multOut[18]), .B1(n16420), .C1(addOut[18]), 
          .D1(addIn2_28__N_1441[18]), .CIN(n18415), .COUT(n18416), .S0(n121[17]), 
          .S1(n121[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_19.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_19.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_19.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_19.INJECT1_1 = "NO";
    PFUMX mux_137_i13 (.BLUT(n588[12]), .ALUT(intgOut3[12]), .C0(n21420), 
          .Z(n618[12])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    CCU2D add_1212_11 (.A0(n5451), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n5453), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18235), 
          .COUT(n18236), .S0(n2373[9]), .S1(n2373[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(126[13] 142[6])
    defparam add_1212_11.INIT0 = 16'hf555;
    defparam add_1212_11.INIT1 = 16'hf555;
    defparam add_1212_11.INJECT1_0 = "NO";
    defparam add_1212_11.INJECT1_1 = "NO";
    CCU2D addOut_2126_add_4_17 (.A0(multOut[15]), .B0(n16420), .C0(addOut[15]), 
          .D0(addIn2_28__N_1441[15]), .A1(multOut[16]), .B1(n16420), .C1(addOut[16]), 
          .D1(addIn2_28__N_1441[16]), .CIN(n18414), .COUT(n18415), .S0(n121[15]), 
          .S1(n121[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126_add_4_17.INIT0 = 16'h569a;
    defparam addOut_2126_add_4_17.INIT1 = 16'h569a;
    defparam addOut_2126_add_4_17.INJECT1_0 = "NO";
    defparam addOut_2126_add_4_17.INJECT1_1 = "NO";
    FD1S3AX addOut_2126__i1 (.D(n121[1]), .CK(clk_N_875), .Q(addOut[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i1.GSR = "ENABLED";
    PFUMX i17351 (.BLUT(n21504), .ALUT(n21505), .C0(n21467), .Z(n16496));
    PFUMX mux_137_i14 (.BLUT(n588[13]), .ALUT(intgOut3[13]), .C0(n21420), 
          .Z(n618[13])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i15 (.BLUT(n588[14]), .ALUT(intgOut3[14]), .C0(n21420), 
          .Z(n618[14])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i16 (.BLUT(n588[15]), .ALUT(intgOut3[15]), .C0(n21420), 
          .Z(n618[15])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i17 (.BLUT(n588[16]), .ALUT(intgOut3[16]), .C0(n21420), 
          .Z(n618[16])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i18 (.BLUT(n588[17]), .ALUT(intgOut3[17]), .C0(n21420), 
          .Z(n618[17])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i19 (.BLUT(n588[18]), .ALUT(intgOut3[18]), .C0(n21420), 
          .Z(n618[18])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i20 (.BLUT(n588[19]), .ALUT(intgOut3[19]), .C0(n21420), 
          .Z(n618[19])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    PFUMX mux_137_i21 (.BLUT(n588[20]), .ALUT(intgOut3[20]), .C0(n21420), 
          .Z(n618[20])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=317, LSE_RLINE=317 */ ;
    FD1S3AX addOut_2126__i2 (.D(n121[2]), .CK(clk_N_875), .Q(addOut[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i2.GSR = "ENABLED";
    FD1S3AX addOut_2126__i3 (.D(n121[3]), .CK(clk_N_875), .Q(addOut[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i3.GSR = "ENABLED";
    FD1S3AX addOut_2126__i4 (.D(n121[4]), .CK(clk_N_875), .Q(addOut[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i4.GSR = "ENABLED";
    FD1S3AX addOut_2126__i5 (.D(n121[5]), .CK(clk_N_875), .Q(addOut[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i5.GSR = "ENABLED";
    FD1S3AX addOut_2126__i6 (.D(n121[6]), .CK(clk_N_875), .Q(addOut[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i6.GSR = "ENABLED";
    FD1S3AX addOut_2126__i7 (.D(n121[7]), .CK(clk_N_875), .Q(addOut[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i7.GSR = "ENABLED";
    FD1S3AX addOut_2126__i8 (.D(n121[8]), .CK(clk_N_875), .Q(addOut[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i8.GSR = "ENABLED";
    FD1S3AX addOut_2126__i9 (.D(n121[9]), .CK(clk_N_875), .Q(addOut[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i9.GSR = "ENABLED";
    FD1S3AX addOut_2126__i10 (.D(n121[10]), .CK(clk_N_875), .Q(addOut[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i10.GSR = "ENABLED";
    FD1S3AX addOut_2126__i11 (.D(n121[11]), .CK(clk_N_875), .Q(addOut[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i11.GSR = "ENABLED";
    FD1S3AX addOut_2126__i12 (.D(n121[12]), .CK(clk_N_875), .Q(addOut[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i12.GSR = "ENABLED";
    FD1S3AX addOut_2126__i13 (.D(n121[13]), .CK(clk_N_875), .Q(addOut[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i13.GSR = "ENABLED";
    FD1S3AX addOut_2126__i14 (.D(n121[14]), .CK(clk_N_875), .Q(addOut[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i14.GSR = "ENABLED";
    FD1S3AX addOut_2126__i15 (.D(n121[15]), .CK(clk_N_875), .Q(addOut[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i15.GSR = "ENABLED";
    FD1S3AX addOut_2126__i16 (.D(n121[16]), .CK(clk_N_875), .Q(addOut[16])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i16.GSR = "ENABLED";
    FD1S3AX addOut_2126__i17 (.D(n121[17]), .CK(clk_N_875), .Q(addOut[17])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i17.GSR = "ENABLED";
    FD1S3AX addOut_2126__i18 (.D(n121[18]), .CK(clk_N_875), .Q(addOut[18])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i18.GSR = "ENABLED";
    FD1S3AX addOut_2126__i19 (.D(n121[19]), .CK(clk_N_875), .Q(addOut[19])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i19.GSR = "ENABLED";
    FD1S3AX addOut_2126__i20 (.D(n121[20]), .CK(clk_N_875), .Q(addOut[20])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i20.GSR = "ENABLED";
    FD1S3AX addOut_2126__i21 (.D(n121[21]), .CK(clk_N_875), .Q(addOut[21])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i21.GSR = "ENABLED";
    FD1S3AX addOut_2126__i22 (.D(n121[22]), .CK(clk_N_875), .Q(addOut[22])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i22.GSR = "ENABLED";
    FD1S3AX addOut_2126__i23 (.D(n121[23]), .CK(clk_N_875), .Q(addOut[23])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i23.GSR = "ENABLED";
    FD1S3AX addOut_2126__i24 (.D(n121[24]), .CK(clk_N_875), .Q(addOut[24])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i24.GSR = "ENABLED";
    FD1S3AX addOut_2126__i25 (.D(n121[25]), .CK(clk_N_875), .Q(addOut[25])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i25.GSR = "ENABLED";
    FD1S3AX addOut_2126__i26 (.D(n121[26]), .CK(clk_N_875), .Q(addOut[26])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i26.GSR = "ENABLED";
    FD1S3AX addOut_2126__i27 (.D(n121[27]), .CK(clk_N_875), .Q(addOut[27])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i27.GSR = "ENABLED";
    FD1S3AX addOut_2126__i28 (.D(n121[28]), .CK(clk_N_875), .Q(addOut[28])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pid.vhd(230[13:19])
    defparam addOut_2126__i28.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWMGENERATOR
//

module PWMGENERATOR (pwm_clk, PWM_m4, LED4_c, clkout_c_enable_362, PWMdut_m4, 
            GND_net);
    input pwm_clk;
    output PWM_m4;
    output LED4_c;
    input clkout_c_enable_362;
    input [9:0]PWMdut_m4;
    input GND_net;
    
    wire pwm_clk /* synthesis SET_AS_NETWORK=pwm_clk, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(88[9:16])
    wire [9:0]cnt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(41[10:13])
    
    wire n14213;
    wire [9:0]n45;
    
    wire PWM_N_2176, free_N_2188, n17, n16, n3892, n11553, n14, 
        n10, n7;
    wire [9:0]n1;
    
    wire n7_adj_2326, n8, n18391, n18390, n18389, n18388, n18387, 
        n21437, n18353, n18352, n18351, n18350, n18349;
    
    FD1S3IX cnt_2130__i0 (.D(n45[0]), .CK(pwm_clk), .CD(n14213), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i0.GSR = "ENABLED";
    FD1S3AX PWM_22 (.D(PWM_N_2176), .CK(pwm_clk), .Q(PWM_m4)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=13, LSE_RCOL=25, LSE_LLINE=358, LSE_RLINE=358 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam PWM_22.GSR = "ENABLED";
    FD1P3AX free_21 (.D(free_N_2188), .SP(clkout_c_enable_362), .CK(pwm_clk), 
            .Q(LED4_c));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(52[2] 80[9])
    defparam free_21.GSR = "DISABLED";
    LUT4 i17189_4_lut (.A(n17), .B(cnt[7]), .C(n16), .D(cnt[3]), .Z(n14213)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(77[6:16])
    defparam i17189_4_lut.init = 16'h0400;
    LUT4 i7_4_lut (.A(cnt[2]), .B(cnt[9]), .C(cnt[5]), .D(cnt[6]), .Z(n17)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    LUT4 i6_4_lut (.A(cnt[1]), .B(cnt[4]), .C(cnt[8]), .D(cnt[0]), .Z(n16)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i6_4_lut.init = 16'hffef;
    LUT4 i1810_1_lut (.A(n3892), .Z(PWM_N_2176)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1810_1_lut.init = 16'h5555;
    LUT4 i6_4_lut_adj_40 (.A(PWMdut_m4[9]), .B(PWMdut_m4[3]), .C(PWMdut_m4[4]), 
         .D(n11553), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i6_4_lut_adj_40.init = 16'hfffe;
    LUT4 i2_2_lut (.A(PWMdut_m4[6]), .B(PWMdut_m4[7]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(PWMdut_m4[2]), .B(PWMdut_m4[1]), .C(PWMdut_m4[0]), 
         .Z(n11553)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i13320_2_lut (.A(PWMdut_m4[8]), .B(n7), .Z(n1[8])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13320_2_lut.init = 16'heeee;
    LUT4 i5_4_lut (.A(PWMdut_m4[9]), .B(n7_adj_2326), .C(PWMdut_m4[7]), 
         .D(n8), .Z(n7)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(PWMdut_m4[6]), .B(n11553), .C(PWMdut_m4[4]), .D(PWMdut_m4[3]), 
         .Z(n7_adj_2326)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut.init = 16'ha8a0;
    LUT4 i2_2_lut_adj_41 (.A(PWMdut_m4[5]), .B(PWMdut_m4[8]), .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_41.init = 16'h8888;
    LUT4 i13318_2_lut (.A(PWMdut_m4[6]), .B(n7), .Z(n1[6])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13318_2_lut.init = 16'heeee;
    LUT4 i13316_2_lut (.A(PWMdut_m4[3]), .B(n7), .Z(n1[3])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(59[4] 63[11])
    defparam i13316_2_lut.init = 16'heeee;
    CCU2D cnt_2130_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18391), .S0(n45[9]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2130_add_4_11.INIT1 = 16'h0000;
    defparam cnt_2130_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2130_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_2130_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18390), 
          .COUT(n18391), .S0(n45[7]), .S1(n45[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2130_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2130_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2130_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_2130_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18389), 
          .COUT(n18390), .S0(n45[5]), .S1(n45[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2130_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2130_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2130_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_2130_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18388), 
          .COUT(n18389), .S0(n45[3]), .S1(n45[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2130_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2130_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2130_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2130_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18387), 
          .COUT(n18388), .S0(n45[1]), .S1(n45[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2130_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2130_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2130_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2130_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n18387), .S1(n45[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2130_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2130_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2130_add_4_1.INJECT1_1 = "NO";
    LUT4 i7_4_lut_rep_336 (.A(PWMdut_m4[5]), .B(n14), .C(n10), .D(PWMdut_m4[8]), 
         .Z(n21437)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam i7_4_lut_rep_336.init = 16'hfffe;
    LUT4 DutyCycle_9__I_0_i20_1_lut_4_lut (.A(PWMdut_m4[5]), .B(n14), .C(n10), 
         .D(PWMdut_m4[8]), .Z(free_N_2188)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(54[6:19])
    defparam DutyCycle_9__I_0_i20_1_lut_4_lut.init = 16'h0001;
    CCU2D sub_1808_add_2_11 (.A0(PWMdut_m4[9]), .B0(n21437), .C0(cnt[9]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18353), .S1(n3892));
    defparam sub_1808_add_2_11.INIT0 = 16'h8787;
    defparam sub_1808_add_2_11.INIT1 = 16'h0000;
    defparam sub_1808_add_2_11.INJECT1_0 = "NO";
    defparam sub_1808_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_9 (.A0(PWMdut_m4[7]), .B0(n21437), .C0(cnt[7]), 
          .D0(GND_net), .A1(n1[8]), .B1(n21437), .C1(cnt[8]), .D1(GND_net), 
          .CIN(n18352), .COUT(n18353));
    defparam sub_1808_add_2_9.INIT0 = 16'h8787;
    defparam sub_1808_add_2_9.INIT1 = 16'h8787;
    defparam sub_1808_add_2_9.INJECT1_0 = "NO";
    defparam sub_1808_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_7 (.A0(PWMdut_m4[5]), .B0(n21437), .C0(cnt[5]), 
          .D0(GND_net), .A1(n1[6]), .B1(n21437), .C1(cnt[6]), .D1(GND_net), 
          .CIN(n18351), .COUT(n18352));
    defparam sub_1808_add_2_7.INIT0 = 16'h8787;
    defparam sub_1808_add_2_7.INIT1 = 16'h8787;
    defparam sub_1808_add_2_7.INJECT1_0 = "NO";
    defparam sub_1808_add_2_7.INJECT1_1 = "NO";
    FD1S3IX cnt_2130__i1 (.D(n45[1]), .CK(pwm_clk), .CD(n14213), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i1.GSR = "ENABLED";
    FD1S3IX cnt_2130__i2 (.D(n45[2]), .CK(pwm_clk), .CD(n14213), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i2.GSR = "ENABLED";
    FD1S3IX cnt_2130__i3 (.D(n45[3]), .CK(pwm_clk), .CD(n14213), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i3.GSR = "ENABLED";
    FD1S3IX cnt_2130__i4 (.D(n45[4]), .CK(pwm_clk), .CD(n14213), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i4.GSR = "ENABLED";
    FD1S3IX cnt_2130__i5 (.D(n45[5]), .CK(pwm_clk), .CD(n14213), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i5.GSR = "ENABLED";
    FD1S3IX cnt_2130__i6 (.D(n45[6]), .CK(pwm_clk), .CD(n14213), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i6.GSR = "ENABLED";
    FD1S3IX cnt_2130__i7 (.D(n45[7]), .CK(pwm_clk), .CD(n14213), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i7.GSR = "ENABLED";
    FD1S3IX cnt_2130__i8 (.D(n45[8]), .CK(pwm_clk), .CD(n14213), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i8.GSR = "ENABLED";
    FD1S3IX cnt_2130__i9 (.D(n45[9]), .CK(pwm_clk), .CD(n14213), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/pwm_gen.vhd(76[9:12])
    defparam cnt_2130__i9.GSR = "ENABLED";
    CCU2D sub_1808_add_2_5 (.A0(n1[3]), .B0(n21437), .C0(cnt[3]), .D0(GND_net), 
          .A1(cnt[4]), .B1(n21437), .C1(n7), .D1(PWMdut_m4[4]), .CIN(n18350), 
          .COUT(n18351));
    defparam sub_1808_add_2_5.INIT0 = 16'h8787;
    defparam sub_1808_add_2_5.INIT1 = 16'h5955;
    defparam sub_1808_add_2_5.INJECT1_0 = "NO";
    defparam sub_1808_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_3 (.A0(cnt[1]), .B0(n21437), .C0(n7), .D0(PWMdut_m4[1]), 
          .A1(cnt[2]), .B1(n21437), .C1(n7), .D1(PWMdut_m4[2]), .CIN(n18349), 
          .COUT(n18350));
    defparam sub_1808_add_2_3.INIT0 = 16'h5955;
    defparam sub_1808_add_2_3.INIT1 = 16'h5955;
    defparam sub_1808_add_2_3.INJECT1_0 = "NO";
    defparam sub_1808_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1808_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(n21437), .C1(n7), .D1(PWMdut_m4[0]), 
          .COUT(n18349));
    defparam sub_1808_add_2_1.INIT0 = 16'h0000;
    defparam sub_1808_add_2_1.INIT1 = 16'h5955;
    defparam sub_1808_add_2_1.INJECT1_0 = "NO";
    defparam sub_1808_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module HALL
//

module HALL (clk_1mhz, \speed_m4[0] , hallsense_m4, clkout_c_enable_266, 
            clkout_c_enable_362, H_A_m4_c, H_B_m4_c, H_C_m4_c, \speed_m4[1] , 
            \speed_m4[2] , \speed_m4[3] , \speed_m4[4] , \speed_m4[5] , 
            \speed_m4[6] , \speed_m4[7] , \speed_m4[8] , \speed_m4[9] , 
            \speed_m4[10] , \speed_m4[11] , \speed_m4[12] , \speed_m4[13] , 
            \speed_m4[14] , \speed_m4[15] , \speed_m4[16] , \speed_m4[17] , 
            \speed_m4[18] , \speed_m4[19] , GND_net, n22206);
    input clk_1mhz;
    output \speed_m4[0] ;
    output [2:0]hallsense_m4;
    input clkout_c_enable_266;
    input clkout_c_enable_362;
    input H_A_m4_c;
    input H_B_m4_c;
    input H_C_m4_c;
    output \speed_m4[1] ;
    output \speed_m4[2] ;
    output \speed_m4[3] ;
    output \speed_m4[4] ;
    output \speed_m4[5] ;
    output \speed_m4[6] ;
    output \speed_m4[7] ;
    output \speed_m4[8] ;
    output \speed_m4[9] ;
    output \speed_m4[10] ;
    output \speed_m4[11] ;
    output \speed_m4[12] ;
    output \speed_m4[13] ;
    output \speed_m4[14] ;
    output \speed_m4[15] ;
    output \speed_m4[16] ;
    output \speed_m4[17] ;
    output \speed_m4[18] ;
    output \speed_m4[19] ;
    input GND_net;
    input n22206;
    
    wire clk_1mhz /* synthesis SET_AS_NETWORK=clk_1mhz, is_clock=1 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/toplevelfinal.vhd(86[9:17])
    wire [6:0]stable_count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(62[10:22])
    
    wire stable_counting, n14464, n21497;
    wire [19:0]speedt;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(61[10:16])
    
    wire clk_1mhz_enable_88;
    wire [19:0]count_19__N_2069;
    
    wire n21496;
    wire [6:0]n63;
    
    wire n21468, n21447;
    wire [19:0]count;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(60[10:15])
    
    wire n4633;
    wire [19:0]speedt_19__N_2049;
    
    wire hall3_lat, n4, n11560, n11568, hall3_old, hall1_lat, hall2_lat, 
        hall1_old, hall2_old, n21417, n21469, stable_counting_N_2131, 
        n4_adj_2324, n19651, n21413, n13, n12, n19879, n19883, 
        n19881, n19715, n21428, n19585, n21429, n18856, n19785, 
        clk_1mhz_enable_187, n25, n26, n22, n19805, n19803, n24, 
        n18, n18323, n18322, n18321, n18320, n18319, n18318, n18317, 
        n18316, n18315, n18314;
    
    FD1P3IX stable_count__i0 (.D(n21497), .SP(stable_counting), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_count[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i0.GSR = "ENABLED";
    FD1P3AX speedt_i0_i0 (.D(count_19__N_2069[0]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i0.GSR = "ENABLED";
    LUT4 i2559_2_lut_rep_395 (.A(stable_count[1]), .B(stable_count[0]), 
         .Z(n21496)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2559_2_lut_rep_395.init = 16'h8888;
    LUT4 i2564_2_lut_3_lut (.A(stable_count[1]), .B(stable_count[0]), .C(stable_count[2]), 
         .Z(n63[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2564_2_lut_3_lut.init = 16'h7878;
    LUT4 i2571_2_lut_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n63[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2571_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2566_2_lut_rep_367_3_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[2]), .Z(n21468)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2566_2_lut_rep_367_3_lut.init = 16'h8080;
    LUT4 i2573_2_lut_rep_346_3_lut_4_lut (.A(stable_count[1]), .B(stable_count[0]), 
         .C(stable_count[3]), .D(stable_count[2]), .Z(n21447)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2573_2_lut_rep_346_3_lut_4_lut.init = 16'h8000;
    FD1S3IX count__i0 (.D(count_19__N_2069[0]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX speed__i1 (.D(speedt_19__N_2049[0]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[0] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i0 (.D(hall3_lat), .CK(clk_1mhz), .Q(hallsense_m4[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i0.GSR = "ENABLED";
    LUT4 i2555_1_lut_rep_396 (.A(stable_count[0]), .Z(n21497)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2555_1_lut_rep_396.init = 16'h5555;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(stable_count[0]), .B(stable_count[4]), 
         .C(n21468), .D(stable_count[3]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D))))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h7ddd;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[0]), 
         .D(speedt[0]), .Z(speedt_19__N_2049[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX hall3_old_56 (.D(hall3_lat), .SP(clkout_c_enable_266), .CK(clk_1mhz), 
            .Q(hall3_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_old_56.GSR = "DISABLED";
    LUT4 mux_9_i2_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[1]), 
         .D(speedt[1]), .Z(speedt_19__N_2049[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[2]), 
         .D(speedt[2]), .Z(speedt_19__N_2049[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[3]), 
         .D(speedt[3]), .Z(speedt_19__N_2049[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[4]), 
         .D(speedt[4]), .Z(speedt_19__N_2049[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[5]), 
         .D(speedt[5]), .Z(speedt_19__N_2049[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[6]), 
         .D(speedt[6]), .Z(speedt_19__N_2049[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[7]), 
         .D(speedt[7]), .Z(speedt_19__N_2049[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i9_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[8]), 
         .D(speedt[8]), .Z(speedt_19__N_2049[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i9_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX hall1_lat_57 (.D(H_A_m4_c), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall1_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_lat_57.GSR = "DISABLED";
    LUT4 mux_9_i10_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[9]), 
         .D(speedt[9]), .Z(speedt_19__N_2049[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i11_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[10]), 
         .D(speedt[10]), .Z(speedt_19__N_2049[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i12_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[11]), 
         .D(speedt[11]), .Z(speedt_19__N_2049[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i12_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX hall2_lat_58 (.D(H_B_m4_c), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall2_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_lat_58.GSR = "DISABLED";
    FD1P3AX hall3_lat_59 (.D(H_C_m4_c), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall3_lat));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall3_lat_59.GSR = "DISABLED";
    LUT4 mux_9_i13_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[12]), 
         .D(speedt[12]), .Z(speedt_19__N_2049[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i13_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX hall1_old_54 (.D(hall1_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall1_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall1_old_54.GSR = "DISABLED";
    LUT4 mux_9_i14_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[13]), 
         .D(speedt[13]), .Z(speedt_19__N_2049[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i15_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[14]), 
         .D(speedt[14]), .Z(speedt_19__N_2049[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i15_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX hall2_old_55 (.D(hall2_lat), .SP(clkout_c_enable_362), .CK(clk_1mhz), 
            .Q(hall2_old));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam hall2_old_55.GSR = "DISABLED";
    LUT4 mux_9_i16_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[15]), 
         .D(speedt[15]), .Z(speedt_19__N_2049[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i17_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[16]), 
         .D(speedt[16]), .Z(speedt_19__N_2049[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i18_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[17]), 
         .D(speedt[17]), .Z(speedt_19__N_2049[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i19_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[18]), 
         .D(speedt[18]), .Z(speedt_19__N_2049[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i20_3_lut_4_lut (.A(n11560), .B(n11568), .C(count_19__N_2069[19]), 
         .D(speedt[19]), .Z(speedt_19__N_2049[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_9_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2585_2_lut_rep_316_3_lut_4_lut (.A(stable_count[3]), .B(n21468), 
         .C(stable_count[5]), .D(stable_count[4]), .Z(n21417)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2585_2_lut_rep_316_3_lut_4_lut.init = 16'h78f0;
    LUT4 i16409_3_lut (.A(n21469), .B(stable_counting), .C(stable_counting_N_2131), 
         .Z(n14464)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16409_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut (.A(hall2_old), .B(hall1_old), .C(hall2_lat), .D(hall1_lat), 
         .Z(n4_adj_2324)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i1_4_lut_adj_37 (.A(n63[2]), .B(n19651), .C(n21413), .D(n4), 
         .Z(stable_counting_N_2131)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(106[7:23])
    defparam i1_4_lut_adj_37.init = 16'h0004;
    LUT4 i2557_2_lut (.A(stable_count[1]), .B(stable_count[0]), .Z(n63[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2557_2_lut.init = 16'h6666;
    LUT4 i11563_4_lut (.A(n11560), .B(n11568), .C(stable_counting), .D(stable_counting_N_2131), 
         .Z(clk_1mhz_enable_88)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C))) */ ;
    defparam i11563_4_lut.init = 16'hcaea;
    LUT4 i7_4_lut (.A(n13), .B(count[8]), .C(n12), .D(count[0]), .Z(n11560)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i5_4_lut (.A(count[9]), .B(count[3]), .C(count[2]), .D(count[13]), 
         .Z(n13)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5_4_lut.init = 16'h8000;
    LUT4 i4_4_lut (.A(count[10]), .B(n19879), .C(n19883), .D(n19881), 
         .Z(n12)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h0002;
    LUT4 i16427_4_lut (.A(count[6]), .B(count[1]), .C(count[7]), .D(n19715), 
         .Z(n19879)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16427_4_lut.init = 16'hfffe;
    LUT4 i16431_4_lut (.A(count[15]), .B(count[19]), .C(count[5]), .D(count[16]), 
         .Z(n19883)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16431_4_lut.init = 16'hfffe;
    LUT4 i16429_4_lut (.A(count[12]), .B(count[4]), .C(count[17]), .D(count[18]), 
         .Z(n19881)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16429_4_lut.init = 16'hfffe;
    LUT4 i16264_2_lut (.A(count[11]), .B(count[14]), .Z(n19715)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16264_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(n19651), .B(stable_count[0]), .C(n21428), .D(n19585), 
         .Z(n11568)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    FD1P3AX speedt_i0_i1 (.D(count_19__N_2069[1]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i1.GSR = "ENABLED";
    FD1P3AX speedt_i0_i2 (.D(count_19__N_2069[2]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i2.GSR = "ENABLED";
    FD1P3AX speedt_i0_i3 (.D(count_19__N_2069[3]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i3.GSR = "ENABLED";
    FD1P3AX speedt_i0_i4 (.D(count_19__N_2069[4]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i4.GSR = "ENABLED";
    FD1P3AX speedt_i0_i5 (.D(count_19__N_2069[5]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i5.GSR = "ENABLED";
    FD1P3AX speedt_i0_i6 (.D(count_19__N_2069[6]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i6.GSR = "ENABLED";
    FD1P3AX speedt_i0_i7 (.D(count_19__N_2069[7]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i7.GSR = "ENABLED";
    FD1P3AX speedt_i0_i8 (.D(count_19__N_2069[8]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i8.GSR = "ENABLED";
    FD1P3AX speedt_i0_i9 (.D(count_19__N_2069[9]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i9.GSR = "ENABLED";
    FD1P3AX speedt_i0_i10 (.D(count_19__N_2069[10]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i10.GSR = "ENABLED";
    FD1P3AX speedt_i0_i11 (.D(count_19__N_2069[11]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i11.GSR = "ENABLED";
    FD1P3AX speedt_i0_i12 (.D(count_19__N_2069[12]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i12.GSR = "ENABLED";
    FD1P3AX speedt_i0_i13 (.D(count_19__N_2069[13]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i13.GSR = "ENABLED";
    FD1P3AX speedt_i0_i14 (.D(count_19__N_2069[14]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i14.GSR = "ENABLED";
    FD1P3AX speedt_i0_i15 (.D(count_19__N_2069[15]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i15.GSR = "ENABLED";
    FD1P3AX speedt_i0_i16 (.D(count_19__N_2069[16]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i16.GSR = "ENABLED";
    FD1P3AX speedt_i0_i17 (.D(count_19__N_2069[17]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i17.GSR = "ENABLED";
    FD1P3AX speedt_i0_i18 (.D(count_19__N_2069[18]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i18.GSR = "ENABLED";
    FD1P3AX speedt_i0_i19 (.D(count_19__N_2069[19]), .SP(clk_1mhz_enable_88), 
            .CK(clk_1mhz), .Q(speedt[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speedt_i0_i19.GSR = "ENABLED";
    LUT4 i2299_2_lut (.A(stable_counting), .B(stable_counting_N_2131), .Z(n4633)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i2299_2_lut.init = 16'h8888;
    FD1S3IX count__i1 (.D(count_19__N_2069[1]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(count_19__N_2069[2]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(count_19__N_2069[3]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(count_19__N_2069[4]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(count_19__N_2069[5]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(count_19__N_2069[6]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(count_19__N_2069[7]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(count_19__N_2069[8]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(count_19__N_2069[9]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(count_19__N_2069[10]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_19__N_2069[11]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(count_19__N_2069[12]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(count_19__N_2069[13]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(count_19__N_2069[14]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(count_19__N_2069[15]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i15.GSR = "ENABLED";
    FD1S3IX count__i16 (.D(count_19__N_2069[16]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i16.GSR = "ENABLED";
    FD1S3IX count__i17 (.D(count_19__N_2069[17]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i17.GSR = "ENABLED";
    FD1S3IX count__i18 (.D(count_19__N_2069[18]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i18.GSR = "ENABLED";
    FD1S3IX count__i19 (.D(count_19__N_2069[19]), .CK(clk_1mhz), .CD(n4633), 
            .Q(count[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam count__i19.GSR = "ENABLED";
    FD1P3AX speed__i2 (.D(speedt_19__N_2049[1]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[1] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i2.GSR = "ENABLED";
    FD1P3AX speed__i3 (.D(speedt_19__N_2049[2]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[2] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i3.GSR = "ENABLED";
    FD1P3AX speed__i4 (.D(speedt_19__N_2049[3]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[3] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i4.GSR = "ENABLED";
    FD1P3AX speed__i5 (.D(speedt_19__N_2049[4]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i5.GSR = "ENABLED";
    FD1P3AX speed__i6 (.D(speedt_19__N_2049[5]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i6.GSR = "ENABLED";
    FD1P3AX speed__i7 (.D(speedt_19__N_2049[6]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i7.GSR = "ENABLED";
    FD1P3AX speed__i8 (.D(speedt_19__N_2049[7]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i8.GSR = "ENABLED";
    FD1P3AX speed__i9 (.D(speedt_19__N_2049[8]), .SP(stable_counting), .CK(clk_1mhz), 
            .Q(\speed_m4[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i9.GSR = "ENABLED";
    FD1P3AX speed__i10 (.D(speedt_19__N_2049[9]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i10.GSR = "ENABLED";
    FD1P3AX speed__i11 (.D(speedt_19__N_2049[10]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i11.GSR = "ENABLED";
    FD1P3AX speed__i12 (.D(speedt_19__N_2049[11]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i12.GSR = "ENABLED";
    FD1P3AX speed__i13 (.D(speedt_19__N_2049[12]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i13.GSR = "ENABLED";
    FD1P3AX speed__i14 (.D(speedt_19__N_2049[13]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i14.GSR = "ENABLED";
    FD1P3AX speed__i15 (.D(speedt_19__N_2049[14]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i15.GSR = "ENABLED";
    FD1P3AX speed__i16 (.D(speedt_19__N_2049[15]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i16.GSR = "ENABLED";
    FD1P3AX speed__i17 (.D(speedt_19__N_2049[16]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i17.GSR = "ENABLED";
    FD1P3AX speed__i18 (.D(speedt_19__N_2049[17]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i18.GSR = "ENABLED";
    FD1P3AX speed__i19 (.D(speedt_19__N_2049[18]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i19.GSR = "ENABLED";
    FD1P3AX speed__i20 (.D(speedt_19__N_2049[19]), .SP(stable_counting), 
            .CK(clk_1mhz), .Q(\speed_m4[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam speed__i20.GSR = "ENABLED";
    FD1S3AY Hall_sns_i1 (.D(hall2_lat), .CK(clk_1mhz), .Q(hallsense_m4[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i1.GSR = "ENABLED";
    FD1S3AY Hall_sns_i2 (.D(hall1_lat), .CK(clk_1mhz), .Q(hallsense_m4[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam Hall_sns_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut (.A(n63[3]), .B(n63[6]), .C(n21417), .D(n63[2]), 
         .Z(n19585)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_312_4_lut (.A(stable_count[5]), .B(n21429), .C(n63[6]), 
         .D(n63[3]), .Z(n21413)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2_3_lut_rep_312_4_lut.init = 16'hfff6;
    LUT4 i17266_4_lut (.A(n18856), .B(n19785), .C(hall3_old), .D(hall3_lat), 
         .Z(clk_1mhz_enable_187)) /* synthesis lut_function=((B+!(C (D)+!C !(D)))+!A) */ ;
    defparam i17266_4_lut.init = 16'hdffd;
    LUT4 i1_4_lut_adj_38 (.A(n25), .B(count[0]), .C(n26), .D(count[10]), 
         .Z(n18856)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i1_4_lut_adj_38.init = 16'hfbff;
    LUT4 i16334_4_lut (.A(hall1_old), .B(hall2_old), .C(hall1_lat), .D(hall2_lat), 
         .Z(n19785)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i16334_4_lut.init = 16'h7bde;
    LUT4 i11_4_lut (.A(count[18]), .B(n22), .C(n19805), .D(n19803), 
         .Z(n25)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i11_4_lut.init = 16'hefff;
    LUT4 i12_4_lut (.A(count[5]), .B(n24), .C(n18), .D(count[19]), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(count[17]), .B(count[16]), .C(count[14]), .D(count[15]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i16353_2_lut (.A(count[8]), .B(count[13]), .Z(n19805)) /* synthesis lut_function=(A (B)) */ ;
    defparam i16353_2_lut.init = 16'h8888;
    LUT4 i16351_3_lut (.A(count[2]), .B(count[3]), .C(count[9]), .Z(n19803)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16351_3_lut.init = 16'h8080;
    LUT4 i10_4_lut (.A(count[11]), .B(count[7]), .C(count[6]), .D(count[1]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i4_2_lut (.A(count[4]), .B(count[12]), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i2578_2_lut_rep_327_3_lut_4_lut (.A(stable_count[2]), .B(n21496), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21428)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2578_2_lut_rep_327_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2580_2_lut_rep_328_3_lut_4_lut (.A(stable_count[2]), .B(n21496), 
         .C(stable_count[4]), .D(stable_count[3]), .Z(n21429)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2580_2_lut_rep_328_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_rep_368 (.A(hall3_old), .B(n4_adj_2324), .C(hall3_lat), 
         .Z(n21469)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i2_3_lut_rep_368.init = 16'hdede;
    LUT4 i1_2_lut_4_lut_adj_39 (.A(hall3_old), .B(n4_adj_2324), .C(hall3_lat), 
         .D(n63[1]), .Z(n19651)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_39.init = 16'h2100;
    LUT4 i2592_3_lut_4_lut (.A(stable_count[4]), .B(n21447), .C(stable_count[5]), 
         .D(stable_count[6]), .Z(n63[6])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(100[21:33])
    defparam i2592_3_lut_4_lut.init = 16'h7f80;
    CCU2D add_7_21 (.A0(count[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18323), 
          .S0(count_19__N_2069[19]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_21.INIT0 = 16'h5aaa;
    defparam add_7_21.INIT1 = 16'h0000;
    defparam add_7_21.INJECT1_0 = "NO";
    defparam add_7_21.INJECT1_1 = "NO";
    CCU2D add_7_19 (.A0(count[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18322), .COUT(n18323), .S0(count_19__N_2069[17]), .S1(count_19__N_2069[18]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_19.INIT0 = 16'h5aaa;
    defparam add_7_19.INIT1 = 16'h5aaa;
    defparam add_7_19.INJECT1_0 = "NO";
    defparam add_7_19.INJECT1_1 = "NO";
    CCU2D add_7_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18321), .COUT(n18322), .S0(count_19__N_2069[15]), .S1(count_19__N_2069[16]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h5aaa;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18320), .COUT(n18321), .S0(count_19__N_2069[13]), .S1(count_19__N_2069[14]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18319), .COUT(n18320), .S0(count_19__N_2069[11]), .S1(count_19__N_2069[12]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18318), .COUT(n18319), .S0(count_19__N_2069[9]), .S1(count_19__N_2069[10]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18317), 
          .COUT(n18318), .S0(count_19__N_2069[7]), .S1(count_19__N_2069[8]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18316), 
          .COUT(n18317), .S0(count_19__N_2069[5]), .S1(count_19__N_2069[6]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18315), 
          .COUT(n18316), .S0(count_19__N_2069[3]), .S1(count_19__N_2069[4]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n18314), 
          .COUT(n18315), .S0(count_19__N_2069[1]), .S1(count_19__N_2069[2]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n18314), 
          .S1(count_19__N_2069[0]));   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(86[12:17])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    FD1P3IX stable_count__i6 (.D(n63[6]), .SP(stable_counting), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_count[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i6.GSR = "ENABLED";
    FD1P3IX stable_count__i5 (.D(n21417), .SP(stable_counting), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_count[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i5.GSR = "ENABLED";
    FD1P3IX stable_count__i4 (.D(n21428), .SP(stable_counting), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_count[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i4.GSR = "ENABLED";
    FD1P3IX stable_count__i3 (.D(n63[3]), .SP(stable_counting), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_count[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i3.GSR = "ENABLED";
    FD1P3IX stable_count__i2 (.D(n63[2]), .SP(stable_counting), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_count[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i2.GSR = "ENABLED";
    FD1P3IX stable_count__i1 (.D(n63[1]), .SP(stable_counting), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_count[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_count__i1.GSR = "ENABLED";
    FD1P3IX stable_counting_62 (.D(n22206), .SP(clk_1mhz_enable_187), .CD(n14464), 
            .CK(clk_1mhz), .Q(stable_counting)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=14, LSE_RCOL=18, LSE_LLINE=352, LSE_RLINE=352 */ ;   // c:/users/gebruiker/workspace/lattice/motorcontroller-prototype/hallinput.vhd(75[2] 121[9])
    defparam stable_counting_62.GSR = "ENABLED";
    
endmodule
